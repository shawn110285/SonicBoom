module Queue_5_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 34016:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 34017:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 34018:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 34019:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34022:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34023:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 34024:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 34025:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 34026:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 34027:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 34028:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 34029:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 34032:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 34047:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 34053:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 34056:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_param_MPORT_data = 2'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_sink_MPORT_data = 1'h0;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_denied_MPORT_data = 1'h0;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 34062:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 34060:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34072:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34071:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34070:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34069:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34068:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34067:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34066:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 34065:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 34021:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34022:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34022:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 34035:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 34048:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34023:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 34023:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 34050:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 34054:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 34024:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 34024:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 34057:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 34058:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 39472:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 39473:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 39474:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [31:0] io_enq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [31:0] io_deq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 39475:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [31:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [31:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [31:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39478:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39479:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39480:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 39481:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 39482:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 39483:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 39484:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39485:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39488:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39503:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39509:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 39512:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_param_MPORT_data = 3'h0;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_source_MPORT_data = 1'h0;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
  assign ram_corrupt_MPORT_data = 1'h0;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 39518:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 39516:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39528:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39527:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39526:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39525:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39524:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39523:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39522:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39521:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39477:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39478:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39478:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 39491:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39504:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39479:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39479:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 39506:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39510:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39480:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39480:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 39513:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 39514:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_7_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 39536:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 39537:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 39538:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [1:0]  io_enq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [3:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [2:0]  io_enq_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [1:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [3:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [2:0]  io_deq_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 39539:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [1:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [1:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [1:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [3:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [3:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [3:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [2:0] ram_sink [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [2:0] ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_sink_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  ram_denied [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_denied_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39542:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39543:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39544:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 39545:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 39546:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 39547:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 39548:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39549:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 39552:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39567:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 39573:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 39576:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sink_io_deq_bits_MPORT_addr = value_1;
  assign ram_sink_io_deq_bits_MPORT_data = ram_sink[ram_sink_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_sink_MPORT_data = io_enq_bits_sink;
  assign ram_sink_MPORT_addr = value;
  assign ram_sink_MPORT_mask = 1'h1;
  assign ram_sink_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_denied_io_deq_bits_MPORT_addr = value_1;
  assign ram_denied_io_deq_bits_MPORT_data = ram_denied[ram_denied_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_denied_MPORT_data = io_enq_bits_denied;
  assign ram_denied_MPORT_addr = value;
  assign ram_denied_MPORT_mask = 1'h1;
  assign ram_denied_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 39582:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 39580:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39592:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39591:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39590:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39589:4]
  assign io_deq_bits_sink = ram_sink_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39588:4]
  assign io_deq_bits_denied = ram_denied_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39587:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39586:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 39585:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_sink_MPORT_en & ram_sink_MPORT_mask) begin
      ram_sink[ram_sink_MPORT_addr] <= ram_sink_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_denied_MPORT_en & ram_denied_MPORT_mask) begin
      ram_denied[ram_denied_MPORT_addr] <= ram_denied_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 39541:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39542:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39542:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 39555:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39568:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39543:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 39543:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 39570:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 39574:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39544:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 39544:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 39577:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 39578:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_denied[initvar] = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HellaPeekingArbiter_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 369217:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 369218:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 369219:4]
  output        io_in_1_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input         io_in_1_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [2:0]  io_in_1_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [2:0]  io_in_1_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [3:0]  io_in_1_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [3:0]  io_in_1_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [63:0] io_in_1_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input         io_in_1_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [7:0]  io_in_1_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input         io_in_1_bits_last, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output        io_in_4_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input         io_in_4_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [2:0]  io_in_4_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [2:0]  io_in_4_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [3:0]  io_in_4_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [3:0]  io_in_4_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [31:0] io_in_4_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [63:0] io_in_4_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input         io_in_4_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input  [7:0]  io_in_4_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input         io_in_4_bits_last, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  input         io_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output        io_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [3:0]  io_out_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [63:0] io_out_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output [7:0]  io_out_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
  output        io_out_bits_last // @[chipyard.TestHarness.SmallBoomConfig.fir 369220:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] lockIdx; // @[Arbiters.scala 25:20 chipyard.TestHarness.SmallBoomConfig.fir 369225:4]
  reg  locked; // @[Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369226:4]
  wire [2:0] choice = io_in_1_valid ? 3'h1 : 3'h4; // @[Mux.scala 47:69 chipyard.TestHarness.SmallBoomConfig.fir 369229:4]
  wire [2:0] chosen = locked ? lockIdx : choice; // @[Arbiters.scala 36:19 chipyard.TestHarness.SmallBoomConfig.fir 369231:4]
  wire  _io_in_1_ready_T = chosen == 3'h1; // @[Arbiters.scala 39:46 chipyard.TestHarness.SmallBoomConfig.fir 369235:4]
  wire  _io_in_4_ready_T = chosen == 3'h4; // @[Arbiters.scala 39:46 chipyard.TestHarness.SmallBoomConfig.fir 369244:4]
  wire [2:0] _GEN_14 = 3'h1 == chosen ? 3'h3 : 3'h4; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_15 = 3'h1 == chosen ? io_in_1_bits_opcode : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_16 = 3'h1 == chosen ? io_in_1_bits_param : 3'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [3:0] _GEN_17 = 3'h1 == chosen ? io_in_1_bits_size : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [3:0] _GEN_18 = 3'h1 == chosen ? io_in_1_bits_source : 4'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [63:0] _GEN_20 = 3'h1 == chosen ? io_in_1_bits_data : 64'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [7:0] _GEN_22 = 3'h1 == chosen ? io_in_1_bits_union : 8'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire  _GEN_23 = 3'h1 == chosen ? io_in_1_bits_last : 1'h1; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire  _GEN_25 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_valid; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_26 = 3'h2 == chosen ? 3'h2 : _GEN_14; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_27 = 3'h2 == chosen ? 3'h0 : _GEN_15; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_28 = 3'h2 == chosen ? 3'h0 : _GEN_16; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [3:0] _GEN_29 = 3'h2 == chosen ? 4'h0 : _GEN_17; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [3:0] _GEN_30 = 3'h2 == chosen ? 4'h0 : _GEN_18; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [63:0] _GEN_32 = 3'h2 == chosen ? 64'h0 : _GEN_20; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire  _GEN_33 = 3'h2 == chosen ? 1'h0 : 3'h1 == chosen & io_in_1_bits_corrupt; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [7:0] _GEN_34 = 3'h2 == chosen ? 8'h0 : _GEN_22; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire  _GEN_37 = 3'h3 == chosen ? 1'h0 : _GEN_25; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_38 = 3'h3 == chosen ? 3'h1 : _GEN_26; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_39 = 3'h3 == chosen ? 3'h0 : _GEN_27; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [2:0] _GEN_40 = 3'h3 == chosen ? 3'h0 : _GEN_28; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [3:0] _GEN_41 = 3'h3 == chosen ? 4'h0 : _GEN_29; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [3:0] _GEN_42 = 3'h3 == chosen ? 4'h0 : _GEN_30; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [63:0] _GEN_44 = 3'h3 == chosen ? 64'h0 : _GEN_32; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire  _GEN_45 = 3'h3 == chosen ? 1'h0 : _GEN_33; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire [7:0] _GEN_46 = 3'h3 == chosen ? 8'h0 : _GEN_34; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369249:4]
  wire  _T_1 = ~locked; // @[Arbiters.scala 59:11 chipyard.TestHarness.SmallBoomConfig.fir 369251:6]
  wire  _GEN_61 = _T_1 | locked; // @[Arbiters.scala 59:50 chipyard.TestHarness.SmallBoomConfig.fir 369253:6 Arbiters.scala 61:14 chipyard.TestHarness.SmallBoomConfig.fir 369255:8 Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369226:4]
  assign io_in_1_ready = io_out_ready & _io_in_1_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.SmallBoomConfig.fir 369236:4]
  assign io_in_4_ready = io_out_ready & _io_in_4_ready_T; // @[Arbiters.scala 39:36 chipyard.TestHarness.SmallBoomConfig.fir 369245:4]
  assign io_out_valid = 3'h4 == chosen ? io_in_4_valid : _GEN_37; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_chanId = 3'h4 == chosen ? 3'h0 : _GEN_38; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_opcode = 3'h4 == chosen ? io_in_4_bits_opcode : _GEN_39; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_param = 3'h4 == chosen ? io_in_4_bits_param : _GEN_40; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_size = 3'h4 == chosen ? io_in_4_bits_size : _GEN_41; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_source = 3'h4 == chosen ? io_in_4_bits_source : _GEN_42; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_address = 3'h4 == chosen ? io_in_4_bits_address : 32'h0; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_data = 3'h4 == chosen ? io_in_4_bits_data : _GEN_44; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_corrupt = 3'h4 == chosen ? io_in_4_bits_corrupt : _GEN_45; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_union = 3'h4 == chosen ? io_in_4_bits_union : _GEN_46; // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  assign io_out_bits_last = 3'h4 == chosen ? io_in_4_bits_last : 3'h3 == chosen | (3'h2 == chosen | _GEN_23); // @[Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4 Arbiters.scala 42:16 chipyard.TestHarness.SmallBoomConfig.fir 369247:4]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiters.scala 25:20 chipyard.TestHarness.SmallBoomConfig.fir 369225:4]
      lockIdx <= 3'h0; // @[Arbiters.scala 25:20 chipyard.TestHarness.SmallBoomConfig.fir 369225:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.SmallBoomConfig.fir 369250:4]
      if (_T_1) begin // @[Arbiters.scala 59:50 chipyard.TestHarness.SmallBoomConfig.fir 369253:6]
        if (io_in_1_valid) begin // @[Mux.scala 47:69 chipyard.TestHarness.SmallBoomConfig.fir 369229:4]
          lockIdx <= 3'h1;
        end else begin
          lockIdx <= 3'h4;
        end
      end
    end
    if (reset) begin // @[Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369226:4]
      locked <= 1'h0; // @[Arbiters.scala 26:19 chipyard.TestHarness.SmallBoomConfig.fir 369226:4]
    end else if (_T) begin // @[Arbiters.scala 58:24 chipyard.TestHarness.SmallBoomConfig.fir 369250:4]
      if (io_out_bits_last) begin // @[Arbiters.scala 64:35 chipyard.TestHarness.SmallBoomConfig.fir 369257:6]
        locked <= 1'h0; // @[Arbiters.scala 65:14 chipyard.TestHarness.SmallBoomConfig.fir 369258:8]
      end else begin
        locked <= _GEN_61;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockIdx = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  locked = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericSerializer_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 369262:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 369263:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 369264:4]
  output        io_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input         io_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [2:0]  io_in_bits_chanId, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [2:0]  io_in_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [2:0]  io_in_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [3:0]  io_in_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [3:0]  io_in_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [31:0] io_in_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [63:0] io_in_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input         io_in_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input  [7:0]  io_in_bits_union, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input         io_in_bits_last, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  input         io_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  output        io_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
  output [3:0]  io_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 369265:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [122:0] data; // @[Serdes.scala 175:17 chipyard.TestHarness.SmallBoomConfig.fir 369267:4]
  reg  sending; // @[Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369268:4]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369269:4]
  reg [4:0] sendCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369270:4]
  wire  wrap_wrap = sendCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 369274:6]
  wire [4:0] _wrap_value_T_1 = sendCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 369276:6]
  wire  sendDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369273:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 369281:6 chipyard.TestHarness.SmallBoomConfig.fir 369272:4]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369288:4]
  wire [122:0] _data_T = {io_in_bits_chanId,io_in_bits_opcode,io_in_bits_param,io_in_bits_size,io_in_bits_source,
    io_in_bits_address,io_in_bits_data,io_in_bits_corrupt,io_in_bits_union,io_in_bits_last}; // @[Serdes.scala 185:24 chipyard.TestHarness.SmallBoomConfig.fir 369298:6]
  wire  _GEN_4 = _T_1 | sending; // @[Serdes.scala 184:23 chipyard.TestHarness.SmallBoomConfig.fir 369289:4 Serdes.scala 186:13 chipyard.TestHarness.SmallBoomConfig.fir 369300:6 Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369268:4]
  wire [122:0] _data_T_1 = {{4'd0}, data[122:4]}; // @[Serdes.scala 189:39 chipyard.TestHarness.SmallBoomConfig.fir 369304:6]
  assign io_in_ready = ~sending; // @[Serdes.scala 180:18 chipyard.TestHarness.SmallBoomConfig.fir 369283:4]
  assign io_out_valid = sending; // @[Serdes.scala 181:16 chipyard.TestHarness.SmallBoomConfig.fir 369285:4]
  assign io_out_bits = data[3:0]; // @[Serdes.scala 182:22 chipyard.TestHarness.SmallBoomConfig.fir 369286:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 189:24 chipyard.TestHarness.SmallBoomConfig.fir 369303:4]
      data <= _data_T_1; // @[Serdes.scala 189:31 chipyard.TestHarness.SmallBoomConfig.fir 369305:6]
    end else if (_T_1) begin // @[Serdes.scala 184:23 chipyard.TestHarness.SmallBoomConfig.fir 369289:4]
      data <= _data_T; // @[Serdes.scala 185:10 chipyard.TestHarness.SmallBoomConfig.fir 369299:6]
    end
    if (reset) begin // @[Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369268:4]
      sending <= 1'h0; // @[Serdes.scala 177:24 chipyard.TestHarness.SmallBoomConfig.fir 369268:4]
    end else if (sendDone) begin // @[Serdes.scala 191:19 chipyard.TestHarness.SmallBoomConfig.fir 369307:4]
      sending <= 1'h0; // @[Serdes.scala 191:29 chipyard.TestHarness.SmallBoomConfig.fir 369308:6]
    end else begin
      sending <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369270:4]
      sendCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369270:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369273:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 369278:6]
        sendCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 369279:8]
      end else begin
        sendCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 369277:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  data = _RAND_0[122:0];
  _RAND_1 = {1{`RANDOM}};
  sending = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericDeserializer_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 369311:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 369312:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 369313:4]
  output        io_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  input         io_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  input  [3:0]  io_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  input         io_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output        io_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [2:0]  io_out_bits_chanId, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [2:0]  io_out_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [2:0]  io_out_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [3:0]  io_out_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [3:0]  io_out_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [31:0] io_out_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [63:0] io_out_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output        io_out_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
  output [7:0]  io_out_bits_union // @[chipyard.TestHarness.SmallBoomConfig.fir 369314:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] data_0; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_1; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_2; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_3; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_4; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_5; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_6; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_7; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_8; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_9; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_10; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_11; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_12; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_13; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_14; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_15; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_16; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_17; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_18; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_19; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_20; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_21; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_22; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_23; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_24; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_25; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_26; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_27; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_28; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_29; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg [3:0] data_30; // @[Serdes.scala 202:17 chipyard.TestHarness.SmallBoomConfig.fir 369316:4]
  reg  receiving; // @[Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369317:4]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369318:4]
  reg [4:0] recvCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369319:4]
  wire  wrap_wrap = recvCount == 5'h1e; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 369323:6]
  wire [4:0] _wrap_value_T_1 = recvCount + 5'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 369325:6]
  wire  recvDone = _T & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369322:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 369330:6 chipyard.TestHarness.SmallBoomConfig.fir 369321:4]
  wire [27:0] io_out_bits_lo_lo = {data_6,data_5,data_4,data_3,data_2,data_1,data_0}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369340:4]
  wire [59:0] io_out_bits_lo = {data_14,data_13,data_12,data_11,data_10,data_9,data_8,data_7,io_out_bits_lo_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369348:4]
  wire [31:0] io_out_bits_hi_lo = {data_22,data_21,data_20,data_19,data_18,data_17,data_16,data_15}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369355:4]
  wire [123:0] _io_out_bits_T = {data_30,data_29,data_28,data_27,data_26,data_25,data_24,data_23,io_out_bits_hi_lo,
    io_out_bits_lo}; // @[Serdes.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 369364:4]
  wire  _GEN_65 = recvDone ? 1'h0 : receiving; // @[Serdes.scala 215:19 chipyard.TestHarness.SmallBoomConfig.fir 369402:4 Serdes.scala 215:31 chipyard.TestHarness.SmallBoomConfig.fir 369403:6 Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369317:4]
  wire  _T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 369405:4]
  wire  _GEN_66 = _T_2 | _GEN_65; // @[Serdes.scala 217:24 chipyard.TestHarness.SmallBoomConfig.fir 369406:4 Serdes.scala 217:36 chipyard.TestHarness.SmallBoomConfig.fir 369407:6]
  assign io_in_ready = receiving; // @[Serdes.scala 207:15 chipyard.TestHarness.SmallBoomConfig.fir 369332:4]
  assign io_out_valid = ~receiving; // @[Serdes.scala 208:19 chipyard.TestHarness.SmallBoomConfig.fir 369333:4]
  assign io_out_bits_chanId = _io_out_bits_T[122:120]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369386:4]
  assign io_out_bits_opcode = _io_out_bits_T[119:117]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369384:4]
  assign io_out_bits_param = _io_out_bits_T[116:114]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369382:4]
  assign io_out_bits_size = _io_out_bits_T[113:110]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369380:4]
  assign io_out_bits_source = _io_out_bits_T[109:106]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369378:4]
  assign io_out_bits_address = _io_out_bits_T[105:74]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369376:4]
  assign io_out_bits_data = _io_out_bits_T[73:10]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369374:4]
  assign io_out_bits_corrupt = _io_out_bits_T[9]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369372:4]
  assign io_out_bits_union = _io_out_bits_T[8:1]; // @[Serdes.scala 209:38 chipyard.TestHarness.SmallBoomConfig.fir 369370:4]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h0 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_0 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h1 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_1 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h2 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_2 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h3 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_3 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h4 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_4 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h5 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_5 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h6 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_6 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h7 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_7 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h8 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_8 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h9 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_9 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'ha == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_10 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'hb == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_11 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'hc == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_12 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'hd == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_13 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'he == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_14 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'hf == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_15 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h10 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_16 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h11 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_17 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h12 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_18 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h13 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_19 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h14 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_20 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h15 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_21 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h16 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_22 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h17 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_23 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h18 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_24 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h19 == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_25 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h1a == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_26 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h1b == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_27 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h1c == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_28 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h1d == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_29 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    if (_T) begin // @[Serdes.scala 211:23 chipyard.TestHarness.SmallBoomConfig.fir 369399:4]
      if (5'h1e == recvCount) begin // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
        data_30 <= io_in_bits; // @[Serdes.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 369400:6]
      end
    end
    receiving <= reset | _GEN_66; // @[Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369317:4 Serdes.scala 204:26 chipyard.TestHarness.SmallBoomConfig.fir 369317:4]
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369319:4]
      recvCount <= 5'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 369319:4]
    end else if (_T) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 369322:4]
      if (wrap_wrap) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 369327:6]
        recvCount <= 5'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 369328:8]
      end else begin
        recvCount <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 369326:6]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  data_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  data_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  data_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  data_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  data_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  data_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  data_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  data_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  data_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  data_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  data_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  data_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  data_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  data_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  data_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  data_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  data_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  data_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  data_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  data_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  data_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  data_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  data_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  data_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  data_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  data_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  data_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  data_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  data_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  data_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  receiving = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  recvCount = _RAND_32[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule



module SerialAdapter_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 380387:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 380388:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 380389:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 380390:4]
  output        io_serial_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380391:4]
  input         io_serial_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380391:4]
  input  [31:0] io_serial_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 380391:4]
  input         io_serial_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 380391:4]
  output        io_serial_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 380391:4]
  output [31:0] io_serial_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 380391:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cmd; // @[SerialAdapter.scala 86:16 chipyard.TestHarness.SmallBoomConfig.fir 380400:4]
  reg [63:0] addr; // @[SerialAdapter.scala 87:17 chipyard.TestHarness.SmallBoomConfig.fir 380401:4]
  reg [63:0] len; // @[SerialAdapter.scala 88:16 chipyard.TestHarness.SmallBoomConfig.fir 380402:4]
  reg [31:0] body_0; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380403:4]
  reg [31:0] body_1; // @[SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380403:4]
  reg [1:0] bodyValid; // @[SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380404:4]
  reg  idx; // @[SerialAdapter.scala 91:16 chipyard.TestHarness.SmallBoomConfig.fir 380405:4]
  reg [3:0] state; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380406:4]
  wire  _io_serial_in_ready_T = state == 4'h0; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380407:4]
  wire  _io_serial_in_ready_T_1 = state == 4'h1; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380408:4]
  wire  _io_serial_in_ready_T_2 = state == 4'h2; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380409:4]
  wire  _io_serial_in_ready_T_3 = state == 4'h6; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380410:4]
  wire  _io_serial_in_ready_T_4 = _io_serial_in_ready_T | _io_serial_in_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380411:4]
  wire  _io_serial_in_ready_T_5 = _io_serial_in_ready_T_4 | _io_serial_in_ready_T_2; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380412:4]
  wire  _io_serial_out_valid_T = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.SmallBoomConfig.fir 380415:4]
  wire [28:0] beatAddr = addr[31:3]; // @[SerialAdapter.scala 103:22 chipyard.TestHarness.SmallBoomConfig.fir 380418:4]
  wire [28:0] nextAddr_hi = beatAddr + 29'h1; // @[SerialAdapter.scala 104:31 chipyard.TestHarness.SmallBoomConfig.fir 380420:4]
  wire [31:0] nextAddr = {nextAddr_hi,3'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380421:4]
  wire [3:0] wmask_lo = bodyValid[0] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.SmallBoomConfig.fir 380425:4]
  wire [3:0] wmask_hi = bodyValid[1] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12 chipyard.TestHarness.SmallBoomConfig.fir 380427:4]
  wire [7:0] wmask = {wmask_hi,wmask_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380428:4]
  wire [63:0] _GEN_55 = {{32'd0}, nextAddr}; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.SmallBoomConfig.fir 380429:4]
  wire [63:0] addr_size = _GEN_55 - addr; // @[SerialAdapter.scala 107:28 chipyard.TestHarness.SmallBoomConfig.fir 380430:4]
  wire [63:0] len_size_hi = len + 64'h1; // @[SerialAdapter.scala 108:26 chipyard.TestHarness.SmallBoomConfig.fir 380432:4]
  wire [65:0] len_size = {len_size_hi,2'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380433:4]
  wire [65:0] _GEN_56 = {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 380434:4]
  wire  _raw_size_T = len_size < _GEN_56; // @[SerialAdapter.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 380434:4]
  wire [65:0] raw_size = _raw_size_T ? len_size : {{2'd0}, addr_size}; // @[SerialAdapter.scala 109:21 chipyard.TestHarness.SmallBoomConfig.fir 380435:4]
  wire  _rsize_T = 66'h1 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 380436:4]
  wire [1:0] _rsize_T_1 = _rsize_T ? 2'h0 : 2'h3; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 380437:4]
  wire  _rsize_T_2 = 66'h2 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 380438:4]
  wire [1:0] _rsize_T_3 = _rsize_T_2 ? 2'h1 : _rsize_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 380439:4]
  wire  _rsize_T_4 = 66'h4 == raw_size; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 380440:4]
  wire [1:0] rsize = _rsize_T_4 ? 2'h2 : _rsize_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 380441:4]
  wire [1:0] _pow2size_T_66 = raw_size[0] + raw_size[1]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380508:4]
  wire [1:0] _pow2size_T_68 = raw_size[2] + raw_size[3]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380510:4]
  wire [2:0] _pow2size_T_70 = _pow2size_T_66 + _pow2size_T_68; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380512:4]
  wire [1:0] _pow2size_T_72 = raw_size[4] + raw_size[5]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380514:4]
  wire [1:0] _pow2size_T_74 = raw_size[6] + raw_size[7]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380516:4]
  wire [2:0] _pow2size_T_76 = _pow2size_T_72 + _pow2size_T_74; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380518:4]
  wire [3:0] _pow2size_T_78 = _pow2size_T_70 + _pow2size_T_76; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380520:4]
  wire [1:0] _pow2size_T_80 = raw_size[8] + raw_size[9]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380522:4]
  wire [1:0] _pow2size_T_82 = raw_size[10] + raw_size[11]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380524:4]
  wire [2:0] _pow2size_T_84 = _pow2size_T_80 + _pow2size_T_82; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380526:4]
  wire [1:0] _pow2size_T_86 = raw_size[12] + raw_size[13]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380528:4]
  wire [1:0] _pow2size_T_88 = raw_size[14] + raw_size[15]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380530:4]
  wire [2:0] _pow2size_T_90 = _pow2size_T_86 + _pow2size_T_88; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380532:4]
  wire [3:0] _pow2size_T_92 = _pow2size_T_84 + _pow2size_T_90; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380534:4]
  wire [4:0] _pow2size_T_94 = _pow2size_T_78 + _pow2size_T_92; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380536:4]
  wire [1:0] _pow2size_T_96 = raw_size[16] + raw_size[17]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380538:4]
  wire [1:0] _pow2size_T_98 = raw_size[18] + raw_size[19]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380540:4]
  wire [2:0] _pow2size_T_100 = _pow2size_T_96 + _pow2size_T_98; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380542:4]
  wire [1:0] _pow2size_T_102 = raw_size[20] + raw_size[21]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380544:4]
  wire [1:0] _pow2size_T_104 = raw_size[22] + raw_size[23]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380546:4]
  wire [2:0] _pow2size_T_106 = _pow2size_T_102 + _pow2size_T_104; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380548:4]
  wire [3:0] _pow2size_T_108 = _pow2size_T_100 + _pow2size_T_106; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380550:4]
  wire [1:0] _pow2size_T_110 = raw_size[24] + raw_size[25]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380552:4]
  wire [1:0] _pow2size_T_112 = raw_size[26] + raw_size[27]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380554:4]
  wire [2:0] _pow2size_T_114 = _pow2size_T_110 + _pow2size_T_112; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380556:4]
  wire [1:0] _pow2size_T_116 = raw_size[28] + raw_size[29]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380558:4]
  wire [1:0] _pow2size_T_118 = raw_size[31] + raw_size[32]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380560:4]
  wire [1:0] _GEN_57 = {{1'd0}, raw_size[30]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380562:4]
  wire [2:0] _pow2size_T_120 = _GEN_57 + _pow2size_T_118; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380562:4]
  wire [2:0] _pow2size_T_122 = _pow2size_T_116 + _pow2size_T_120[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380564:4]
  wire [3:0] _pow2size_T_124 = _pow2size_T_114 + _pow2size_T_122; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380566:4]
  wire [4:0] _pow2size_T_126 = _pow2size_T_108 + _pow2size_T_124; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380568:4]
  wire [5:0] _pow2size_T_128 = _pow2size_T_94 + _pow2size_T_126; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380570:4]
  wire [1:0] _pow2size_T_130 = raw_size[33] + raw_size[34]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380572:4]
  wire [1:0] _pow2size_T_132 = raw_size[35] + raw_size[36]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380574:4]
  wire [2:0] _pow2size_T_134 = _pow2size_T_130 + _pow2size_T_132; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380576:4]
  wire [1:0] _pow2size_T_136 = raw_size[37] + raw_size[38]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380578:4]
  wire [1:0] _pow2size_T_138 = raw_size[39] + raw_size[40]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380580:4]
  wire [2:0] _pow2size_T_140 = _pow2size_T_136 + _pow2size_T_138; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380582:4]
  wire [3:0] _pow2size_T_142 = _pow2size_T_134 + _pow2size_T_140; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380584:4]
  wire [1:0] _pow2size_T_144 = raw_size[41] + raw_size[42]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380586:4]
  wire [1:0] _pow2size_T_146 = raw_size[43] + raw_size[44]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380588:4]
  wire [2:0] _pow2size_T_148 = _pow2size_T_144 + _pow2size_T_146; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380590:4]
  wire [1:0] _pow2size_T_150 = raw_size[45] + raw_size[46]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380592:4]
  wire [1:0] _pow2size_T_152 = raw_size[47] + raw_size[48]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380594:4]
  wire [2:0] _pow2size_T_154 = _pow2size_T_150 + _pow2size_T_152; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380596:4]
  wire [3:0] _pow2size_T_156 = _pow2size_T_148 + _pow2size_T_154; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380598:4]
  wire [4:0] _pow2size_T_158 = _pow2size_T_142 + _pow2size_T_156; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380600:4]
  wire [1:0] _pow2size_T_160 = raw_size[49] + raw_size[50]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380602:4]
  wire [1:0] _pow2size_T_162 = raw_size[51] + raw_size[52]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380604:4]
  wire [2:0] _pow2size_T_164 = _pow2size_T_160 + _pow2size_T_162; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380606:4]
  wire [1:0] _pow2size_T_166 = raw_size[53] + raw_size[54]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380608:4]
  wire [1:0] _pow2size_T_168 = raw_size[55] + raw_size[56]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380610:4]
  wire [2:0] _pow2size_T_170 = _pow2size_T_166 + _pow2size_T_168; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380612:4]
  wire [3:0] _pow2size_T_172 = _pow2size_T_164 + _pow2size_T_170; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380614:4]
  wire [1:0] _pow2size_T_174 = raw_size[57] + raw_size[58]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380616:4]
  wire [1:0] _pow2size_T_176 = raw_size[59] + raw_size[60]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380618:4]
  wire [2:0] _pow2size_T_178 = _pow2size_T_174 + _pow2size_T_176; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380620:4]
  wire [1:0] _pow2size_T_180 = raw_size[61] + raw_size[62]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380622:4]
  wire [1:0] _pow2size_T_182 = raw_size[64] + raw_size[65]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380624:4]
  wire [1:0] _GEN_58 = {{1'd0}, raw_size[63]}; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380626:4]
  wire [2:0] _pow2size_T_184 = _GEN_58 + _pow2size_T_182; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380626:4]
  wire [2:0] _pow2size_T_186 = _pow2size_T_180 + _pow2size_T_184[1:0]; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380628:4]
  wire [3:0] _pow2size_T_188 = _pow2size_T_178 + _pow2size_T_186; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380630:4]
  wire [4:0] _pow2size_T_190 = _pow2size_T_172 + _pow2size_T_188; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380632:4]
  wire [5:0] _pow2size_T_192 = _pow2size_T_158 + _pow2size_T_190; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380634:4]
  wire [6:0] _pow2size_T_194 = _pow2size_T_128 + _pow2size_T_192; // @[Bitwise.scala 47:55 chipyard.TestHarness.SmallBoomConfig.fir 380636:4]
  wire  pow2size = _pow2size_T_194 == 7'h1; // @[SerialAdapter.scala 113:37 chipyard.TestHarness.SmallBoomConfig.fir 380638:4]
  wire [2:0] byteAddr = pow2size ? addr[2:0] : 3'h0; // @[SerialAdapter.scala 114:21 chipyard.TestHarness.SmallBoomConfig.fir 380640:4]
  wire [31:0] put_acquire_address = {beatAddr, 3'h0}; // @[SerialAdapter.scala 117:19 chipyard.TestHarness.SmallBoomConfig.fir 380641:4]
  wire [63:0] put_acquire_data = {body_1,body_0}; // @[SerialAdapter.scala 118:10 chipyard.TestHarness.SmallBoomConfig.fir 380642:4]
  wire [31:0] get_acquire_address = {beatAddr,byteAddr}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380707:4]
  wire [2:0] _get_acquire_a_mask_sizeOH_T = {{1'd0}, rsize}; // @[Misc.scala 201:34 chipyard.TestHarness.SmallBoomConfig.fir 380773:4]
  wire [1:0] get_acquire_a_mask_sizeOH_shiftAmount = _get_acquire_a_mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 380774:4]
  wire [3:0] _get_acquire_a_mask_sizeOH_T_1 = 4'h1 << get_acquire_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 380775:4]
  wire [2:0] get_acquire_a_mask_sizeOH = _get_acquire_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 380777:4]
  wire  _get_acquire_a_mask_T = rsize >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 380778:4]
  wire  get_acquire_a_mask_size = get_acquire_a_mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 380779:4]
  wire  get_acquire_a_mask_bit = get_acquire_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 380780:4]
  wire  get_acquire_a_mask_nbit = ~get_acquire_a_mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 380781:4]
  wire  _get_acquire_a_mask_acc_T = get_acquire_a_mask_size & get_acquire_a_mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380783:4]
  wire  get_acquire_a_mask_acc = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380784:4]
  wire  _get_acquire_a_mask_acc_T_1 = get_acquire_a_mask_size & get_acquire_a_mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380786:4]
  wire  get_acquire_a_mask_acc_1 = _get_acquire_a_mask_T | _get_acquire_a_mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380787:4]
  wire  get_acquire_a_mask_size_1 = get_acquire_a_mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 380788:4]
  wire  get_acquire_a_mask_bit_1 = get_acquire_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 380789:4]
  wire  get_acquire_a_mask_nbit_1 = ~get_acquire_a_mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 380790:4]
  wire  get_acquire_a_mask_eq_2 = get_acquire_a_mask_nbit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380791:4]
  wire  _get_acquire_a_mask_acc_T_2 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380792:4]
  wire  get_acquire_a_mask_acc_2 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380793:4]
  wire  get_acquire_a_mask_eq_3 = get_acquire_a_mask_nbit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380794:4]
  wire  _get_acquire_a_mask_acc_T_3 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380795:4]
  wire  get_acquire_a_mask_acc_3 = get_acquire_a_mask_acc | _get_acquire_a_mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380796:4]
  wire  get_acquire_a_mask_eq_4 = get_acquire_a_mask_bit & get_acquire_a_mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380797:4]
  wire  _get_acquire_a_mask_acc_T_4 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380798:4]
  wire  get_acquire_a_mask_acc_4 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380799:4]
  wire  get_acquire_a_mask_eq_5 = get_acquire_a_mask_bit & get_acquire_a_mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380800:4]
  wire  _get_acquire_a_mask_acc_T_5 = get_acquire_a_mask_size_1 & get_acquire_a_mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380801:4]
  wire  get_acquire_a_mask_acc_5 = get_acquire_a_mask_acc_1 | _get_acquire_a_mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380802:4]
  wire  get_acquire_a_mask_size_2 = get_acquire_a_mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 380803:4]
  wire  get_acquire_a_mask_bit_2 = get_acquire_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 380804:4]
  wire  get_acquire_a_mask_nbit_2 = ~get_acquire_a_mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 380805:4]
  wire  get_acquire_a_mask_eq_6 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380806:4]
  wire  _get_acquire_a_mask_acc_T_6 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380807:4]
  wire  get_acquire_a_mask_lo_lo_lo = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380808:4]
  wire  get_acquire_a_mask_eq_7 = get_acquire_a_mask_eq_2 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380809:4]
  wire  _get_acquire_a_mask_acc_T_7 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380810:4]
  wire  get_acquire_a_mask_lo_lo_hi = get_acquire_a_mask_acc_2 | _get_acquire_a_mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380811:4]
  wire  get_acquire_a_mask_eq_8 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380812:4]
  wire  _get_acquire_a_mask_acc_T_8 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380813:4]
  wire  get_acquire_a_mask_lo_hi_lo = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380814:4]
  wire  get_acquire_a_mask_eq_9 = get_acquire_a_mask_eq_3 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380815:4]
  wire  _get_acquire_a_mask_acc_T_9 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380816:4]
  wire  get_acquire_a_mask_lo_hi_hi = get_acquire_a_mask_acc_3 | _get_acquire_a_mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380817:4]
  wire  get_acquire_a_mask_eq_10 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380818:4]
  wire  _get_acquire_a_mask_acc_T_10 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380819:4]
  wire  get_acquire_a_mask_hi_lo_lo = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380820:4]
  wire  get_acquire_a_mask_eq_11 = get_acquire_a_mask_eq_4 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380821:4]
  wire  _get_acquire_a_mask_acc_T_11 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380822:4]
  wire  get_acquire_a_mask_hi_lo_hi = get_acquire_a_mask_acc_4 | _get_acquire_a_mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380823:4]
  wire  get_acquire_a_mask_eq_12 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380824:4]
  wire  _get_acquire_a_mask_acc_T_12 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380825:4]
  wire  get_acquire_a_mask_hi_hi_lo = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380826:4]
  wire  get_acquire_a_mask_eq_13 = get_acquire_a_mask_eq_5 & get_acquire_a_mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 380827:4]
  wire  _get_acquire_a_mask_acc_T_13 = get_acquire_a_mask_size_2 & get_acquire_a_mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 380828:4]
  wire  get_acquire_a_mask_hi_hi_hi = get_acquire_a_mask_acc_5 | _get_acquire_a_mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 380829:4]
  wire [7:0] get_acquire_mask = {get_acquire_a_mask_hi_hi_hi,get_acquire_a_mask_hi_hi_lo,get_acquire_a_mask_hi_lo_hi,
    get_acquire_a_mask_hi_lo_lo,get_acquire_a_mask_lo_hi_hi,get_acquire_a_mask_lo_hi_lo,get_acquire_a_mask_lo_lo_hi,
    get_acquire_a_mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380836:4]
  wire  _bundleOut_0_a_valid_T = state == 4'h7; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380840:4]
  wire  _bundleOut_0_a_valid_T_1 = state == 4'h3; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380841:4]
  wire [3:0] get_acquire_size = {{2'd0}, rsize}; // @[Edges.scala 447:17 chipyard.TestHarness.SmallBoomConfig.fir 380766:4 Edges.scala 450:15 chipyard.TestHarness.SmallBoomConfig.fir 380770:4]
  wire  _bundleOut_0_d_ready_T = state == 4'h8; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380860:4]
  wire  _bundleOut_0_d_ready_T_1 = state == 4'h4; // @[package.scala 15:47 chipyard.TestHarness.SmallBoomConfig.fir 380861:4]
  wire  _T_1 = _io_serial_in_ready_T & io_serial_in_valid; // @[SerialAdapter.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 380868:4]
  wire  _GEN_3 = _T_1 ? 1'h0 : idx; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380869:4 SerialAdapter.scala 140:9 chipyard.TestHarness.SmallBoomConfig.fir 380871:6 SerialAdapter.scala 91:16 chipyard.TestHarness.SmallBoomConfig.fir 380405:4]
  wire [63:0] _GEN_4 = _T_1 ? 64'h0 : addr; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380869:4 SerialAdapter.scala 141:10 chipyard.TestHarness.SmallBoomConfig.fir 380872:6 SerialAdapter.scala 87:17 chipyard.TestHarness.SmallBoomConfig.fir 380401:4]
  wire [63:0] _GEN_5 = _T_1 ? 64'h0 : len; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380869:4 SerialAdapter.scala 142:9 chipyard.TestHarness.SmallBoomConfig.fir 380873:6 SerialAdapter.scala 88:16 chipyard.TestHarness.SmallBoomConfig.fir 380402:4]
  wire [3:0] _GEN_6 = _T_1 ? 4'h1 : state; // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380869:4 SerialAdapter.scala 143:11 chipyard.TestHarness.SmallBoomConfig.fir 380874:6 SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380406:4]
  wire  _T_3 = _io_serial_in_ready_T_1 & io_serial_in_valid; // @[SerialAdapter.scala 146:26 chipyard.TestHarness.SmallBoomConfig.fir 380877:4]
  wire [5:0] _addr_T = {idx,5'h0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 380880:6]
  wire [94:0] _GEN_59 = {{63'd0}, io_serial_in_bits}; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.SmallBoomConfig.fir 380881:6]
  wire [94:0] _addr_T_1 = _GEN_59 << _addr_T; // @[SerialAdapter.scala 132:12 chipyard.TestHarness.SmallBoomConfig.fir 380881:6]
  wire [94:0] _GEN_60 = {{31'd0}, addr}; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 380882:6]
  wire [94:0] _addr_T_2 = _GEN_60 | _addr_T_1; // @[SerialAdapter.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 380882:6]
  wire  _idx_T_1 = idx + 1'h1; // @[SerialAdapter.scala 148:16 chipyard.TestHarness.SmallBoomConfig.fir 380885:6]
  wire  _GEN_7 = idx ? 1'h0 : _idx_T_1; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.SmallBoomConfig.fir 380888:6 SerialAdapter.scala 150:11 chipyard.TestHarness.SmallBoomConfig.fir 380889:8 SerialAdapter.scala 148:9 chipyard.TestHarness.SmallBoomConfig.fir 380886:6]
  wire [3:0] _GEN_8 = idx ? 4'h2 : _GEN_6; // @[SerialAdapter.scala 149:43 chipyard.TestHarness.SmallBoomConfig.fir 380888:6 SerialAdapter.scala 151:13 chipyard.TestHarness.SmallBoomConfig.fir 380890:8]
  wire [94:0] _GEN_9 = _T_3 ? _addr_T_2 : {{31'd0}, _GEN_4}; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.SmallBoomConfig.fir 380878:4 SerialAdapter.scala 147:10 chipyard.TestHarness.SmallBoomConfig.fir 380883:6]
  wire  _GEN_10 = _T_3 ? _GEN_7 : _GEN_3; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.SmallBoomConfig.fir 380878:4]
  wire [3:0] _GEN_11 = _T_3 ? _GEN_8 : _GEN_6; // @[SerialAdapter.scala 146:49 chipyard.TestHarness.SmallBoomConfig.fir 380878:4]
  wire  _T_6 = _io_serial_in_ready_T_2 & io_serial_in_valid; // @[SerialAdapter.scala 155:25 chipyard.TestHarness.SmallBoomConfig.fir 380894:4]
  wire [94:0] _GEN_62 = {{31'd0}, len}; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.SmallBoomConfig.fir 380899:6]
  wire [94:0] _len_T_2 = _GEN_62 | _addr_T_1; // @[SerialAdapter.scala 156:16 chipyard.TestHarness.SmallBoomConfig.fir 380899:6]
  wire  _T_8 = cmd == 32'h1; // @[SerialAdapter.scala 160:17 chipyard.TestHarness.SmallBoomConfig.fir 380908:8]
  wire  _T_9 = cmd == 32'h0; // @[SerialAdapter.scala 163:24 chipyard.TestHarness.SmallBoomConfig.fir 380914:10]
  wire  _T_12 = ~reset; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380921:12]
  wire [3:0] _GEN_12 = _T_9 ? 4'h3 : _GEN_11; // @[SerialAdapter.scala 163:38 chipyard.TestHarness.SmallBoomConfig.fir 380915:10 SerialAdapter.scala 164:15 chipyard.TestHarness.SmallBoomConfig.fir 380916:12]
  wire [1:0] _GEN_13 = _T_8 ? 2'h0 : bodyValid; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.SmallBoomConfig.fir 380909:8 SerialAdapter.scala 161:19 chipyard.TestHarness.SmallBoomConfig.fir 380910:10 SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380404:4]
  wire [3:0] _GEN_14 = _T_8 ? 4'h6 : _GEN_12; // @[SerialAdapter.scala 160:32 chipyard.TestHarness.SmallBoomConfig.fir 380909:8 SerialAdapter.scala 162:15 chipyard.TestHarness.SmallBoomConfig.fir 380911:10]
  wire  _GEN_15 = idx ? addr[2] : _idx_T_1; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.SmallBoomConfig.fir 380905:6 SerialAdapter.scala 159:11 chipyard.TestHarness.SmallBoomConfig.fir 380907:8 SerialAdapter.scala 157:9 chipyard.TestHarness.SmallBoomConfig.fir 380903:6]
  wire [1:0] _GEN_16 = idx ? _GEN_13 : bodyValid; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.SmallBoomConfig.fir 380905:6 SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380404:4]
  wire [3:0] _GEN_17 = idx ? _GEN_14 : _GEN_11; // @[SerialAdapter.scala 158:43 chipyard.TestHarness.SmallBoomConfig.fir 380905:6]
  wire [94:0] _GEN_18 = _T_6 ? _len_T_2 : {{31'd0}, _GEN_5}; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380895:4 SerialAdapter.scala 156:9 chipyard.TestHarness.SmallBoomConfig.fir 380900:6]
  wire  _GEN_19 = _T_6 ? _GEN_15 : _GEN_10; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380895:4]
  wire [1:0] _GEN_20 = _T_6 ? _GEN_16 : bodyValid; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380895:4 SerialAdapter.scala 90:22 chipyard.TestHarness.SmallBoomConfig.fir 380404:4]
  wire [3:0] _GEN_21 = _T_6 ? _GEN_17 : _GEN_11; // @[SerialAdapter.scala 155:48 chipyard.TestHarness.SmallBoomConfig.fir 380895:4]
  wire  _T_14 = _bundleOut_0_a_valid_T_1 & auto_out_a_ready; // @[SerialAdapter.scala 171:30 chipyard.TestHarness.SmallBoomConfig.fir 380930:4]
  wire [3:0] _GEN_22 = _T_14 ? 4'h4 : _GEN_21; // @[SerialAdapter.scala 171:46 chipyard.TestHarness.SmallBoomConfig.fir 380931:4 SerialAdapter.scala 172:11 chipyard.TestHarness.SmallBoomConfig.fir 380932:6]
  wire  _T_16 = _bundleOut_0_d_ready_T_1 & auto_out_d_valid; // @[SerialAdapter.scala 175:31 chipyard.TestHarness.SmallBoomConfig.fir 380935:4]
  wire [31:0] _GEN_23 = _T_16 ? auto_out_d_bits_data[31:0] : body_0; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380936:4 SerialAdapter.scala 176:10 chipyard.TestHarness.SmallBoomConfig.fir 380944:6 SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380403:4]
  wire [31:0] _GEN_24 = _T_16 ? auto_out_d_bits_data[63:32] : body_1; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380936:4 SerialAdapter.scala 176:10 chipyard.TestHarness.SmallBoomConfig.fir 380945:6 SerialAdapter.scala 89:17 chipyard.TestHarness.SmallBoomConfig.fir 380403:4]
  wire  _GEN_25 = _T_16 ? addr[2] : _GEN_19; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380936:4 SerialAdapter.scala 177:9 chipyard.TestHarness.SmallBoomConfig.fir 380947:6]
  wire [94:0] _GEN_26 = _T_16 ? {{63'd0}, nextAddr} : _GEN_9; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380936:4 SerialAdapter.scala 178:10 chipyard.TestHarness.SmallBoomConfig.fir 380948:6]
  wire [3:0] _GEN_27 = _T_16 ? 4'h5 : _GEN_22; // @[SerialAdapter.scala 175:47 chipyard.TestHarness.SmallBoomConfig.fir 380936:4 SerialAdapter.scala 179:11 chipyard.TestHarness.SmallBoomConfig.fir 380949:6]
  wire  _T_20 = _io_serial_out_valid_T & io_serial_out_ready; // @[SerialAdapter.scala 182:31 chipyard.TestHarness.SmallBoomConfig.fir 380952:4]
  wire [63:0] _len_T_4 = len - 64'h1; // @[SerialAdapter.scala 184:16 chipyard.TestHarness.SmallBoomConfig.fir 380958:6]
  wire  _T_21 = len == 64'h0; // @[SerialAdapter.scala 185:15 chipyard.TestHarness.SmallBoomConfig.fir 380960:6]
  wire [3:0] _GEN_28 = idx ? 4'h3 : _GEN_27; // @[SerialAdapter.scala 186:48 chipyard.TestHarness.SmallBoomConfig.fir 380966:8 SerialAdapter.scala 186:56 chipyard.TestHarness.SmallBoomConfig.fir 380967:10]
  wire [3:0] _GEN_29 = _T_21 ? 4'h0 : _GEN_28; // @[SerialAdapter.scala 185:24 chipyard.TestHarness.SmallBoomConfig.fir 380961:6 SerialAdapter.scala 185:32 chipyard.TestHarness.SmallBoomConfig.fir 380962:8]
  wire  _GEN_30 = _T_20 ? _idx_T_1 : _GEN_25; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.SmallBoomConfig.fir 380953:4 SerialAdapter.scala 183:9 chipyard.TestHarness.SmallBoomConfig.fir 380956:6]
  wire [94:0] _GEN_31 = _T_20 ? {{31'd0}, _len_T_4} : _GEN_18; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.SmallBoomConfig.fir 380953:4 SerialAdapter.scala 184:9 chipyard.TestHarness.SmallBoomConfig.fir 380959:6]
  wire [3:0] _GEN_32 = _T_20 ? _GEN_29 : _GEN_27; // @[SerialAdapter.scala 182:55 chipyard.TestHarness.SmallBoomConfig.fir 380953:4]
  wire  _T_24 = _io_serial_in_ready_T_3 & io_serial_in_valid; // @[SerialAdapter.scala 189:32 chipyard.TestHarness.SmallBoomConfig.fir 380971:4]
  wire [1:0] _bodyValid_T = 2'h1 << idx; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 380974:6]
  wire [1:0] _bodyValid_T_1 = bodyValid | _bodyValid_T; // @[SerialAdapter.scala 191:28 chipyard.TestHarness.SmallBoomConfig.fir 380975:6]
  wire  _T_27 = idx | _T_21; // @[SerialAdapter.scala 192:42 chipyard.TestHarness.SmallBoomConfig.fir 380979:6]
  wire [3:0] _GEN_35 = _T_27 ? 4'h7 : _GEN_32; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 380980:6 SerialAdapter.scala 193:13 chipyard.TestHarness.SmallBoomConfig.fir 380981:8]
  wire  _GEN_36 = _T_27 ? _GEN_30 : _idx_T_1; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 380980:6 SerialAdapter.scala 195:11 chipyard.TestHarness.SmallBoomConfig.fir 380986:8]
  wire [94:0] _GEN_37 = _T_27 ? _GEN_31 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 380980:6 SerialAdapter.scala 196:11 chipyard.TestHarness.SmallBoomConfig.fir 380989:8]
  wire [1:0] _GEN_40 = _T_24 ? _bodyValid_T_1 : _GEN_20; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 380972:4 SerialAdapter.scala 191:15 chipyard.TestHarness.SmallBoomConfig.fir 380976:6]
  wire  _GEN_42 = _T_24 ? _GEN_36 : _GEN_30; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 380972:4]
  wire [94:0] _GEN_43 = _T_24 ? _GEN_37 : _GEN_31; // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 380972:4]
  wire  _T_29 = _bundleOut_0_a_valid_T & auto_out_a_ready; // @[SerialAdapter.scala 200:32 chipyard.TestHarness.SmallBoomConfig.fir 380993:4]
  wire  _T_31 = _bundleOut_0_d_ready_T & auto_out_d_valid; // @[SerialAdapter.scala 204:31 chipyard.TestHarness.SmallBoomConfig.fir 380998:4]
  wire [94:0] _GEN_46 = _T_21 ? _GEN_26 : {{63'd0}, nextAddr}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381001:6 SerialAdapter.scala 208:12 chipyard.TestHarness.SmallBoomConfig.fir 381005:8]
  wire [94:0] _GEN_47 = _T_21 ? _GEN_43 : {{31'd0}, _len_T_4}; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381001:6 SerialAdapter.scala 209:11 chipyard.TestHarness.SmallBoomConfig.fir 381008:8]
  wire  _GEN_48 = _T_21 & _GEN_42; // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381001:6 SerialAdapter.scala 210:11 chipyard.TestHarness.SmallBoomConfig.fir 381009:8]
  wire [94:0] _GEN_51 = _T_31 ? _GEN_46 : _GEN_26; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 380999:4]
  wire [94:0] _GEN_52 = _T_31 ? _GEN_47 : _GEN_43; // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 380999:4]
  wire  _GEN_67 = _T_6 & idx & ~_T_8 & ~_T_9; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380923:14]
  assign auto_out_a_valid = _bundleOut_0_a_valid_T | _bundleOut_0_a_valid_T_1; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380842:4]
  assign auto_out_a_bits_opcode = _bundleOut_0_a_valid_T ? 3'h1 : 3'h4; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380845:4]
  assign auto_out_a_bits_size = _bundleOut_0_a_valid_T ? 4'h3 : get_acquire_size; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380845:4]
  assign auto_out_a_bits_address = _bundleOut_0_a_valid_T ? put_acquire_address : get_acquire_address; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380845:4]
  assign auto_out_a_bits_mask = _bundleOut_0_a_valid_T ? wmask : get_acquire_mask; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380845:4]
  assign auto_out_a_bits_data = _bundleOut_0_a_valid_T ? put_acquire_data : 64'h0; // @[SerialAdapter.scala 124:20 chipyard.TestHarness.SmallBoomConfig.fir 380845:4]
  assign auto_out_d_ready = _bundleOut_0_d_ready_T | _bundleOut_0_d_ready_T_1; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380862:4]
  assign io_serial_in_ready = _io_serial_in_ready_T_5 | _io_serial_in_ready_T_3; // @[package.scala 72:59 chipyard.TestHarness.SmallBoomConfig.fir 380413:4]
  assign io_serial_out_valid = state == 4'h5; // @[SerialAdapter.scala 100:32 chipyard.TestHarness.SmallBoomConfig.fir 380415:4]
  assign io_serial_out_bits = idx ? body_1 : body_0; // @[SerialAdapter.scala 101:22 chipyard.TestHarness.SmallBoomConfig.fir 380417:4 SerialAdapter.scala 101:22 chipyard.TestHarness.SmallBoomConfig.fir 380417:4]
  always @(posedge clock) begin
    if (_T_1) begin // @[SerialAdapter.scala 138:48 chipyard.TestHarness.SmallBoomConfig.fir 380869:4]
      cmd <= io_serial_in_bits; // @[SerialAdapter.scala 139:9 chipyard.TestHarness.SmallBoomConfig.fir 380870:6]
    end
    addr <= _GEN_51[63:0];
    len <= _GEN_52[63:0];
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 380972:4]
      if (~idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 380973:6]
        body_0 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 380973:6]
      end else begin
        body_0 <= _GEN_23;
      end
    end else begin
      body_0 <= _GEN_23;
    end
    if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 380972:4]
      if (idx) begin // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 380973:6]
        body_1 <= io_serial_in_bits; // @[SerialAdapter.scala 190:15 chipyard.TestHarness.SmallBoomConfig.fir 380973:6]
      end else begin
        body_1 <= _GEN_24;
      end
    end else begin
      body_1 <= _GEN_24;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 380999:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381001:6]
        bodyValid <= _GEN_40;
      end else begin
        bodyValid <= 2'h0; // @[SerialAdapter.scala 211:17 chipyard.TestHarness.SmallBoomConfig.fir 381010:8]
      end
    end else begin
      bodyValid <= _GEN_40;
    end
    if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 380999:4]
      idx <= _GEN_48;
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 380972:4]
      if (_T_27) begin // @[SerialAdapter.scala 192:58 chipyard.TestHarness.SmallBoomConfig.fir 380980:6]
        idx <= _GEN_30;
      end else begin
        idx <= _idx_T_1; // @[SerialAdapter.scala 195:11 chipyard.TestHarness.SmallBoomConfig.fir 380986:8]
      end
    end else begin
      idx <= _GEN_30;
    end
    if (reset) begin // @[SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380406:4]
      state <= 4'h0; // @[SerialAdapter.scala 97:22 chipyard.TestHarness.SmallBoomConfig.fir 380406:4]
    end else if (_T_31) begin // @[SerialAdapter.scala 204:47 chipyard.TestHarness.SmallBoomConfig.fir 380999:4]
      if (_T_21) begin // @[SerialAdapter.scala 205:24 chipyard.TestHarness.SmallBoomConfig.fir 381001:6]
        state <= 4'h0; // @[SerialAdapter.scala 206:13 chipyard.TestHarness.SmallBoomConfig.fir 381002:8]
      end else begin
        state <= 4'h6; // @[SerialAdapter.scala 212:13 chipyard.TestHarness.SmallBoomConfig.fir 381011:8]
      end
    end else if (_T_29) begin // @[SerialAdapter.scala 200:48 chipyard.TestHarness.SmallBoomConfig.fir 380994:4]
      state <= 4'h8; // @[SerialAdapter.scala 201:11 chipyard.TestHarness.SmallBoomConfig.fir 380995:6]
    end else if (_T_24) begin // @[SerialAdapter.scala 189:55 chipyard.TestHarness.SmallBoomConfig.fir 380972:4]
      state <= _GEN_35;
    end else begin
      state <= _GEN_32;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & idx & ~_T_8 & ~_T_9 & _T_12) begin
          $fwrite(32'h80000002,
            "Assertion failed: Bad TSI command\n    at SerialAdapter.scala:166 assert(false.B, \"Bad TSI command\")\n"); // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380923:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_12) begin
          $fatal; // @[SerialAdapter.scala 166:15 chipyard.TestHarness.SmallBoomConfig.fir 380924:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  len = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  body_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  body_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  bodyValid = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  idx = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_53_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 381031:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 381032:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 381033:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input  [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 381034:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 382973:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 383280:4]
  wire  _source_ok_T = ~io_in_a_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.SmallBoomConfig.fir 381045:6]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 381050:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 381052:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 381053:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 381053:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 381054:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 381056:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 381057:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 381059:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 381060:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 381061:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 381062:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 381063:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381065:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381066:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381068:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381069:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 381070:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 381071:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 381072:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381073:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381074:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381075:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381076:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381077:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381078:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381079:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381080:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381081:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381082:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381083:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381084:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 381085:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 381086:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 381087:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381088:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381089:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381090:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381091:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381092:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381093:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381094:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381095:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381096:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381097:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381098:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381099:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381100:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381101:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381102:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381103:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381104:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381105:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381106:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381107:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381108:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 381109:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 381110:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 381111:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 381118:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381122:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 381134:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 381137:8]
  wire  _T_20 = _T_17 & _source_ok_T; // @[Parameters.scala 1160:30 chipyard.TestHarness.SmallBoomConfig.fir 381140:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381146:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381147:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381148:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381149:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381151:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381152:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381153:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381154:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381156:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381157:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381158:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381159:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381161:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381162:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381163:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381164:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381166:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381167:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381168:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381169:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381171:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381172:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381173:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381174:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381176:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381177:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381178:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.SmallBoomConfig.fir 381185:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381187:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381188:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381190:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381191:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 381192:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 381193:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh10000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 381195:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 381196:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381197:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381198:8]
  wire  _T_81 = _T_20 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.SmallBoomConfig.fir 381201:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381203:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381204:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381271:8]
  wire  _T_149 = _source_ok_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381277:8]
  wire  _T_150 = ~_T_149; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381278:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381285:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381286:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381292:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381293:8]
  wire  _T_158 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 381298:8]
  wire  _T_160 = _T_158 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381300:8]
  wire  _T_161 = ~_T_160; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381301:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 381306:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 381307:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381309:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381310:8]
  wire  _T_167 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 381315:8]
  wire  _T_169 = _T_167 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381317:8]
  wire  _T_170 = ~_T_169; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381318:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 381324:6]
  wire  _T_318 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 381496:8]
  wire  _T_320 = _T_318 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381498:8]
  wire  _T_321 = ~_T_320; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381499:8]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 381522:6]
  wire  _T_339 = _T_20 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381531:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381532:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381546:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 381548:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381591:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381592:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381593:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381594:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381595:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381596:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381597:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381598:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 381600:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381602:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381603:8]
  wire  _T_414 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 381622:8]
  wire  _T_416 = _T_414 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381624:8]
  wire  _T_417 = ~_T_416; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381625:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 381630:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381632:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381633:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 381647:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381704:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381705:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381706:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381707:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381708:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381709:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381710:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 381719:8]
  wire  _T_499 = _T_20 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 381721:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381723:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381724:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 381760:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 381864:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 381865:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 381866:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381868:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381869:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 381875:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 381884:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381928:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381929:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381930:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381931:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381932:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 381933:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 381934:8]
  wire  _T_678 = _T_20 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.SmallBoomConfig.fir 381944:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381946:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381947:8]
  wire  _T_688 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 381966:8]
  wire  _T_690 = _T_688 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381968:8]
  wire  _T_691 = ~_T_690; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381969:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 381983:6]
  wire  _T_774 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 382074:8]
  wire  _T_776 = _T_774 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382076:8]
  wire  _T_777 = ~_T_776; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382077:8]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 382091:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 382161:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 382164:8]
  wire  _T_855 = _T_20 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.SmallBoomConfig.fir 382165:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382167:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382168:8]
  wire  _T_865 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 382187:8]
  wire  _T_867 = _T_865 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382189:8]
  wire  _T_868 = ~_T_867; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382190:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 382214:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382216:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382217:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.SmallBoomConfig.fir 382222:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 382227:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382230:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382231:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 382236:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382238:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382239:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 382244:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382246:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382247:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 382252:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382254:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382255:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 382260:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382262:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382263:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 382269:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 382293:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382295:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382296:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 382301:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382303:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382304:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 382327:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 382368:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382370:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382371:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 382386:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 382421:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 382457:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 382523:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 382528:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 382530:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382532:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382534:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382535:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 382546:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 382547:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 382548:4]
  reg  source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 382549:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 382550:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 382551:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 382552:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 382554:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382556:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382557:6]
  wire  _T_1028 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 382562:6]
  wire  _T_1030 = _T_1028 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382564:6]
  wire  _T_1031 = ~_T_1030; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382565:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 382570:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382572:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382573:6]
  wire  _T_1036 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 382578:6]
  wire  _T_1038 = _T_1036 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382580:6]
  wire  _T_1039 = ~_T_1038; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382581:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 382586:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382588:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382589:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 382596:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 382604:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 382606:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 382608:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 382609:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 382610:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382612:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382614:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382615:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 382626:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 382627:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 382628:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 382629:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 382630:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 382631:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 382632:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 382633:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 382635:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382637:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382638:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 382643:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382645:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382646:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 382651:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382653:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382654:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 382659:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382661:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382662:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 382667:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382669:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382670:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 382675:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382677:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382678:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 382685:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 382694:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 382695:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 382696:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382706:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382708:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382709:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382728:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 382730:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 382731:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 382752:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 382752:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 382753:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 382757:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 382758:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 382758:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 382759:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.SmallBoomConfig.fir 382763:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 382764:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 382768:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 382769:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 382769:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 382770:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 382794:4]
  wire [1:0] _a_set_wo_ready_T = 2'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 382797:6]
  wire [1:0] _GEN_15 = _T_1074 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 382796:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 382798:6 chipyard.TestHarness.SmallBoomConfig.fir 382745:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 382801:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 382806:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 382807:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 382809:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 382810:6]
  wire [2:0] _GEN_77 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 382812:6]
  wire [3:0] _a_opcodes_set_T = {{1'd0}, _GEN_77}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 382812:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382803:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 382808:6 chipyard.TestHarness.SmallBoomConfig.fir 382791:4]
  wire [18:0] _GEN_78 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 382813:6]
  wire [18:0] _a_opcodes_set_T_1 = _GEN_78 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 382813:6]
  wire [3:0] _a_sizes_set_T = {io_in_a_bits_source, 3'h0}; // @[Monitor.scala 657:77 chipyard.TestHarness.SmallBoomConfig.fir 382815:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382803:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 382811:6 chipyard.TestHarness.SmallBoomConfig.fir 382793:4]
  wire [19:0] _GEN_79 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 382816:6]
  wire [19:0] _a_sizes_set_T_1 = _GEN_79 << _a_sizes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 382816:6]
  wire  _T_1079 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 382818:6]
  wire  _T_1081 = ~_T_1079; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 382820:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382822:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382823:6]
  wire [1:0] _GEN_16 = _T_1077 ? _a_set_wo_ready_T : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382803:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 382805:6 chipyard.TestHarness.SmallBoomConfig.fir 382743:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382803:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 382814:6 chipyard.TestHarness.SmallBoomConfig.fir 382747:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 382803:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 382817:6 chipyard.TestHarness.SmallBoomConfig.fir 382749:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 382838:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 382840:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 382841:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 382843:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 382842:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 382844:6 chipyard.TestHarness.SmallBoomConfig.fir 382832:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 382847:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 382850:4]
  wire [30:0] _GEN_81 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 382859:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_81 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 382859:6]
  wire [30:0] _GEN_82 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 382866:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_82 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 382866:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 382851:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 382853:6 chipyard.TestHarness.SmallBoomConfig.fir 382830:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 382851:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 382860:6 chipyard.TestHarness.SmallBoomConfig.fir 382834:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 382851:4 Monitor.scala 678:21 chipyard.TestHarness.SmallBoomConfig.fir 382867:6 chipyard.TestHarness.SmallBoomConfig.fir 382836:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 382876:6]
  wire  same_cycle_resp = _T_1074 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 382877:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 382878:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 382880:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382882:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382883:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 382889:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382890:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382890:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382890:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382890:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 382890:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 382891:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382893:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382894:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 382899:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382901:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382902:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382750:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 382760:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 382910:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382912:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382912:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382912:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382912:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 382912:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 382913:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382915:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382916:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382761:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 382771:4]
  wire [7:0] _GEN_83 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 382921:8]
  wire  _T_1122 = _GEN_83 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 382921:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382923:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382924:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 382932:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 382933:4]
  wire  _T_1130 = _T_1128 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 382935:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 382937:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 382939:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 382940:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382942:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382943:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382744:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382831:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 382949:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 382950:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 382951:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 382952:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382954:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382955:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382742:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 382960:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382829:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 382961:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 382962:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382746:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 382964:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382833:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 382965:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 382966:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382748:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 382968:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 382835:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.SmallBoomConfig.fir 382969:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 382970:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 382972:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 382975:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 382976:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 382977:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 382978:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 382979:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 382980:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382982:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382983:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 382989:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 382993:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 382999:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383034:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 383036:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 383037:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 383070:4]
  wire [15:0] _GEN_87 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 383075:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_87 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 383075:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 383076:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 383154:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 383156:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 383162:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 383164:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 383165:4 Monitor.scala 786:21 chipyard.TestHarness.SmallBoomConfig.fir 383181:6 chipyard.TestHarness.SmallBoomConfig.fir 383152:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 383200:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383204:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383205:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 383058:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 383077:4]
  wire  _T_1194 = _GEN_83 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 383223:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383225:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383226:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 383151:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.SmallBoomConfig.fir 383276:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 383277:4]
  wire  _GEN_93 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381206:10]
  wire  _GEN_109 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381396:10]
  wire  _GEN_127 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381534:10]
  wire  _GEN_141 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381726:10]
  wire  _GEN_151 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381839:10]
  wire  _GEN_161 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381949:10]
  wire  _GEN_171 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382057:10]
  wire  _GEN_181 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382170:10]
  wire  _GEN_193 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382233:10]
  wire  _GEN_203 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382275:10]
  wire  _GEN_213 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382333:10]
  wire  _GEN_223 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382392:10]
  wire  _GEN_229 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382427:10]
  wire  _GEN_235 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382463:10]
  wire  _GEN_241 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382896:10]
  wire  _GEN_246 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382918:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 382973:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 383280:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382532:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382532:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382542:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382543:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382531:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382597:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 382598:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382597:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 382599:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382597:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 382600:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382597:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 382601:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 382597:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 382602:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382612:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382612:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382622:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382623:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382611:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382686:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 382687:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382686:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 382688:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382686:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 382689:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382686:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 382690:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382686:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 382691:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 382686:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 382692:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 382694:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 382694:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 382963:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 382695:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 382695:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 382967:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 382696:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 382696:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 382971:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382706:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382706:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382716:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382717:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382531:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382728:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 382728:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 382738:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 382739:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382611:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 382972:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 382972:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 382994:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 382995:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 382990:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 382999:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 382999:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 383278:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383034:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383034:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 383044:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 383045:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 382611:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381206:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381207:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381273:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381274:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381280:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381281:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381288:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381289:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381295:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381296:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381303:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381304:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381312:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381313:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381320:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_93 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381321:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381396:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381397:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381463:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381464:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381470:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381471:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381478:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381479:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381485:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381486:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381493:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_161) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381494:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381501:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_321) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381502:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381510:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381511:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381518:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_109 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381519:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381534:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381535:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381605:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381606:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381612:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381613:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381619:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381620:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381627:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381628:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381635:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381636:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381643:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_127 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381644:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381726:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381727:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381733:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381734:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381740:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381741:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381748:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381749:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381756:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_141 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381757:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381839:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381840:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381846:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381847:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381853:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381854:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381861:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_417) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381862:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381871:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_151 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381872:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381949:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381950:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381956:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381957:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381963:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381964:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381971:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_691) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381972:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381979:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_161 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 381980:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382057:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382058:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382064:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382065:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382071:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382072:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382079:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_777) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382080:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382087:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_171 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382088:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382170:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382171:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382177:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_150) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382178:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382184:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382185:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382192:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_868) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382193:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382200:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382201:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382208:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_181 & _T_170) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382209:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382219:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382220:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382233:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382234:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382241:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382242:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382249:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382250:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382257:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382258:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382265:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_193 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382266:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382275:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382276:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382290:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382291:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382298:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382299:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382306:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382307:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382314:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382315:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382333:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382334:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382348:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382349:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382356:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382357:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382364:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382365:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382373:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_213 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382374:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382392:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382393:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382400:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382401:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382408:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_223 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382409:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382427:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382428:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382435:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382436:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382444:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_229 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382445:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382463:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382464:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382471:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382472:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382479:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_235 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382480:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382559:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382560:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382567:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1031) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382568:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382575:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382576:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382583:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1039) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382584:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382591:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382592:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382640:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382641:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382648:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382649:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382656:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382657:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382664:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382665:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382672:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382673:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382680:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382681:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382825:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382826:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382885:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382886:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382896:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382897:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382904:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_241 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382905:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382918:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382919:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382926:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_246 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382927:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382945:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382946:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 6 (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382957:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 382958:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382985:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 382986:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383207:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383208:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:25)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383228:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 383229:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inflight_opcodes = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  inflight_sizes = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_20[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerdesser_1_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 383500:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 383501:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 383502:4]
  output        auto_manager_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_manager_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [2:0]  auto_manager_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [2:0]  auto_manager_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [3:0]  auto_manager_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_manager_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [31:0] auto_manager_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [7:0]  auto_manager_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [63:0] auto_manager_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_manager_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_manager_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        auto_manager_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [2:0]  auto_manager_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [1:0]  auto_manager_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [3:0]  auto_manager_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        auto_manager_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [2:0]  auto_manager_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        auto_manager_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [63:0] auto_manager_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        auto_manager_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_client_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        auto_client_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [2:0]  auto_client_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [2:0]  auto_client_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [2:0]  auto_client_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [3:0]  auto_client_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [28:0] auto_client_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [7:0]  auto_client_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output [63:0] auto_client_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        auto_client_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        auto_client_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_client_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [2:0]  auto_client_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [1:0]  auto_client_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [2:0]  auto_client_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [3:0]  auto_client_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_client_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_client_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input  [63:0] auto_client_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  input         auto_client_out_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383503:4]
  output        io_ser_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383504:4]
  input         io_ser_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383504:4]
  input  [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 383504:4]
  input         io_ser_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383504:4]
  output        io_ser_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383504:4]
  output [3:0]  io_ser_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 383504:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
  wire  outArb_clock; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_reset; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_1_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_1_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [2:0] outArb_io_in_1_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [2:0] outArb_io_in_1_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [3:0] outArb_io_in_1_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [3:0] outArb_io_in_1_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [63:0] outArb_io_in_1_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_1_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [7:0] outArb_io_in_1_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_1_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_4_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_4_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [2:0] outArb_io_in_4_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [2:0] outArb_io_in_4_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [3:0] outArb_io_in_4_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [3:0] outArb_io_in_4_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [31:0] outArb_io_in_4_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [63:0] outArb_io_in_4_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_4_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [7:0] outArb_io_in_4_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_in_4_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_out_ready; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_out_valid; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [2:0] outArb_io_out_bits_chanId; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [2:0] outArb_io_out_bits_opcode; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [2:0] outArb_io_out_bits_param; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [3:0] outArb_io_out_bits_size; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [3:0] outArb_io_out_bits_source; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [31:0] outArb_io_out_bits_address; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [63:0] outArb_io_out_bits_data; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_out_bits_corrupt; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire [7:0] outArb_io_out_bits_union; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outArb_io_out_bits_last; // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
  wire  outSer_clock; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  outSer_reset; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  outSer_io_in_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  outSer_io_in_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [2:0] outSer_io_in_bits_chanId; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [2:0] outSer_io_in_bits_opcode; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [2:0] outSer_io_in_bits_param; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [3:0] outSer_io_in_bits_size; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [3:0] outSer_io_in_bits_source; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [31:0] outSer_io_in_bits_address; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [63:0] outSer_io_in_bits_data; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  outSer_io_in_bits_corrupt; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [7:0] outSer_io_in_bits_union; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  outSer_io_in_bits_last; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  outSer_io_out_ready; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  outSer_io_out_valid; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire [3:0] outSer_io_out_bits; // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
  wire  inDes_clock; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire  inDes_reset; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire  inDes_io_in_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire  inDes_io_in_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [3:0] inDes_io_in_bits; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire  inDes_io_out_ready; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire  inDes_io_out_valid; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [2:0] inDes_io_out_bits_chanId; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [2:0] inDes_io_out_bits_opcode; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [2:0] inDes_io_out_bits_param; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [3:0] inDes_io_out_bits_size; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [3:0] inDes_io_out_bits_source; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [31:0] inDes_io_out_bits_address; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [63:0] inDes_io_out_bits_data; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire  inDes_io_out_bits_corrupt; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [7:0] inDes_io_out_bits_union; // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
  wire [1:0] _merged_bits_merged_union_T_1 = {auto_client_out_d_bits_sink,auto_client_out_d_bits_denied}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 383603:4]
  wire  merged_1_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383592:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383788:4]
  wire  _merged_bits_last_T_1 = merged_1_ready & auto_client_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 383616:4]
  wire [12:0] _merged_bits_last_beats1_decode_T_1 = 13'h3f << auto_client_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 383618:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_3 = ~_merged_bits_last_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 383620:4]
  wire [2:0] merged_bits_last_beats1_decode = _merged_bits_last_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 383621:4]
  wire  merged_bits_last_beats1_opdata = auto_client_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 383622:4]
  wire [2:0] merged_bits_last_beats1 = merged_bits_last_beats1_opdata ? merged_bits_last_beats1_decode : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383623:4]
  reg [2:0] merged_bits_last_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383624:4]
  wire [2:0] merged_bits_last_counter1_1 = merged_bits_last_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 383626:4]
  wire  merged_bits_last_first_1 = merged_bits_last_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 383627:4]
  wire  _merged_bits_last_last_T_2 = merged_bits_last_counter_1 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.SmallBoomConfig.fir 383628:4]
  wire  _merged_bits_last_last_T_3 = merged_bits_last_beats1 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.SmallBoomConfig.fir 383629:4]
  wire  merged_4_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383735:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383797:4]
  wire  _merged_bits_last_T_4 = merged_4_ready & auto_manager_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 383758:4]
  wire [20:0] _merged_bits_last_beats1_decode_T_13 = 21'h3f << auto_manager_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 383760:4]
  wire [5:0] _merged_bits_last_beats1_decode_T_15 = ~_merged_bits_last_beats1_decode_T_13[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 383762:4]
  wire [2:0] merged_bits_last_beats1_decode_3 = _merged_bits_last_beats1_decode_T_15[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 383763:4]
  wire  merged_bits_last_beats1_opdata_3 = ~auto_manager_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 383765:4]
  wire [2:0] merged_bits_last_beats1_3 = merged_bits_last_beats1_opdata_3 ? merged_bits_last_beats1_decode_3 : 3'h0; // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383766:4]
  reg [2:0] merged_bits_last_counter_4; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383767:4]
  wire [2:0] merged_bits_last_counter1_4 = merged_bits_last_counter_4 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 383769:4]
  wire  merged_bits_last_first_4 = merged_bits_last_counter_4 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 383770:4]
  wire  _merged_bits_last_last_T_8 = merged_bits_last_counter_4 == 3'h1; // @[Edges.scala 231:25 chipyard.TestHarness.SmallBoomConfig.fir 383771:4]
  wire  _merged_bits_last_last_T_9 = merged_bits_last_beats1_3 == 3'h0; // @[Edges.scala 231:47 chipyard.TestHarness.SmallBoomConfig.fir 383772:4]
  wire  _bundleOut_0_a_valid_T = inDes_io_out_bits_chanId == 3'h0; // @[Serdes.scala 236:37 chipyard.TestHarness.SmallBoomConfig.fir 383810:4]
  wire  _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3; // @[Serdes.scala 239:37 chipyard.TestHarness.SmallBoomConfig.fir 383876:4]
  wire [7:0] _bundleIn_0_d_bits_d_sink_T = {{1'd0}, inDes_io_out_bits_union[7:1]}; // @[Serdes.scala 468:31 chipyard.TestHarness.SmallBoomConfig.fir 383886:4]
  wire  _inDes_io_out_ready_T = 3'h0 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383915:4]
  wire  _inDes_io_out_ready_T_1 = _inDes_io_out_ready_T & auto_client_out_a_ready; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383916:4]
  wire  _inDes_io_out_ready_T_2 = 3'h1 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383917:4]
  wire  _inDes_io_out_ready_T_3 = _inDes_io_out_ready_T_2 ? 1'h0 : _inDes_io_out_ready_T_1; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383918:4]
  wire  _inDes_io_out_ready_T_4 = 3'h2 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383919:4]
  wire  _inDes_io_out_ready_T_5 = _inDes_io_out_ready_T_4 ? 1'h0 : _inDes_io_out_ready_T_3; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383920:4]
  wire  _inDes_io_out_ready_T_6 = 3'h3 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383921:4]
  wire  _inDes_io_out_ready_T_7 = _inDes_io_out_ready_T_6 ? auto_manager_in_d_ready : _inDes_io_out_ready_T_5; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383922:4]
  wire  _inDes_io_out_ready_T_8 = 3'h4 == inDes_io_out_bits_chanId; // @[Mux.scala 80:60 chipyard.TestHarness.SmallBoomConfig.fir 383923:4]
  TLMonitor_53_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 383514:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  HellaPeekingArbiter_inTestHarness outArb ( // @[Serdes.scala 622:24 chipyard.TestHarness.SmallBoomConfig.fir 383545:4]
    .clock(outArb_clock),
    .reset(outArb_reset),
    .io_in_1_ready(outArb_io_in_1_ready),
    .io_in_1_valid(outArb_io_in_1_valid),
    .io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
    .io_in_1_bits_param(outArb_io_in_1_bits_param),
    .io_in_1_bits_size(outArb_io_in_1_bits_size),
    .io_in_1_bits_source(outArb_io_in_1_bits_source),
    .io_in_1_bits_data(outArb_io_in_1_bits_data),
    .io_in_1_bits_corrupt(outArb_io_in_1_bits_corrupt),
    .io_in_1_bits_union(outArb_io_in_1_bits_union),
    .io_in_1_bits_last(outArb_io_in_1_bits_last),
    .io_in_4_ready(outArb_io_in_4_ready),
    .io_in_4_valid(outArb_io_in_4_valid),
    .io_in_4_bits_opcode(outArb_io_in_4_bits_opcode),
    .io_in_4_bits_param(outArb_io_in_4_bits_param),
    .io_in_4_bits_size(outArb_io_in_4_bits_size),
    .io_in_4_bits_source(outArb_io_in_4_bits_source),
    .io_in_4_bits_address(outArb_io_in_4_bits_address),
    .io_in_4_bits_data(outArb_io_in_4_bits_data),
    .io_in_4_bits_corrupt(outArb_io_in_4_bits_corrupt),
    .io_in_4_bits_union(outArb_io_in_4_bits_union),
    .io_in_4_bits_last(outArb_io_in_4_bits_last),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits_chanId(outArb_io_out_bits_chanId),
    .io_out_bits_opcode(outArb_io_out_bits_opcode),
    .io_out_bits_param(outArb_io_out_bits_param),
    .io_out_bits_size(outArb_io_out_bits_size),
    .io_out_bits_source(outArb_io_out_bits_source),
    .io_out_bits_address(outArb_io_out_bits_address),
    .io_out_bits_data(outArb_io_out_bits_data),
    .io_out_bits_corrupt(outArb_io_out_bits_corrupt),
    .io_out_bits_union(outArb_io_out_bits_union),
    .io_out_bits_last(outArb_io_out_bits_last)
  );
  GenericSerializer_inTestHarness outSer ( // @[Serdes.scala 624:24 chipyard.TestHarness.SmallBoomConfig.fir 383548:4]
    .clock(outSer_clock),
    .reset(outSer_reset),
    .io_in_ready(outSer_io_in_ready),
    .io_in_valid(outSer_io_in_valid),
    .io_in_bits_chanId(outSer_io_in_bits_chanId),
    .io_in_bits_opcode(outSer_io_in_bits_opcode),
    .io_in_bits_param(outSer_io_in_bits_param),
    .io_in_bits_size(outSer_io_in_bits_size),
    .io_in_bits_source(outSer_io_in_bits_source),
    .io_in_bits_address(outSer_io_in_bits_address),
    .io_in_bits_data(outSer_io_in_bits_data),
    .io_in_bits_corrupt(outSer_io_in_bits_corrupt),
    .io_in_bits_union(outSer_io_in_bits_union),
    .io_in_bits_last(outSer_io_in_bits_last),
    .io_out_ready(outSer_io_out_ready),
    .io_out_valid(outSer_io_out_valid),
    .io_out_bits(outSer_io_out_bits)
  );
  GenericDeserializer_inTestHarness inDes ( // @[Serdes.scala 629:23 chipyard.TestHarness.SmallBoomConfig.fir 383804:4]
    .clock(inDes_clock),
    .reset(inDes_reset),
    .io_in_ready(inDes_io_in_ready),
    .io_in_valid(inDes_io_in_valid),
    .io_in_bits(inDes_io_in_bits),
    .io_out_ready(inDes_io_out_ready),
    .io_out_valid(inDes_io_out_valid),
    .io_out_bits_chanId(inDes_io_out_bits_chanId),
    .io_out_bits_opcode(inDes_io_out_bits_opcode),
    .io_out_bits_param(inDes_io_out_bits_param),
    .io_out_bits_size(inDes_io_out_bits_size),
    .io_out_bits_source(inDes_io_out_bits_source),
    .io_out_bits_address(inDes_io_out_bits_address),
    .io_out_bits_data(inDes_io_out_bits_data),
    .io_out_bits_corrupt(inDes_io_out_bits_corrupt),
    .io_out_bits_union(inDes_io_out_bits_union)
  );
  assign auto_manager_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383735:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383797:4]
  assign auto_manager_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.SmallBoomConfig.fir 383877:4]
  assign auto_manager_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 461:15 chipyard.TestHarness.SmallBoomConfig.fir 383880:4]
  assign auto_manager_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 462:15 chipyard.TestHarness.SmallBoomConfig.fir 383881:4]
  assign auto_manager_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 463:15 chipyard.TestHarness.SmallBoomConfig.fir 383882:4]
  assign auto_manager_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 464:15 chipyard.TestHarness.SmallBoomConfig.fir 383883:4]
  assign auto_manager_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 468:17 chipyard.TestHarness.SmallBoomConfig.fir 383887:4]
  assign auto_manager_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.SmallBoomConfig.fir 383888:4]
  assign auto_manager_in_d_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 465:15 chipyard.TestHarness.SmallBoomConfig.fir 383884:4]
  assign auto_manager_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 467:17 chipyard.TestHarness.SmallBoomConfig.fir 383885:4]
  assign auto_client_out_a_valid = inDes_io_out_valid & _bundleOut_0_a_valid_T; // @[Serdes.scala 631:45 chipyard.TestHarness.SmallBoomConfig.fir 383811:4]
  assign auto_client_out_a_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 375:15 chipyard.TestHarness.SmallBoomConfig.fir 383814:4]
  assign auto_client_out_a_bits_param = inDes_io_out_bits_param; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 376:15 chipyard.TestHarness.SmallBoomConfig.fir 383815:4]
  assign auto_client_out_a_bits_size = inDes_io_out_bits_size[2:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 377:15 chipyard.TestHarness.SmallBoomConfig.fir 383816:4]
  assign auto_client_out_a_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 378:15 chipyard.TestHarness.SmallBoomConfig.fir 383817:4]
  assign auto_client_out_a_bits_address = inDes_io_out_bits_address[28:0]; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 379:15 chipyard.TestHarness.SmallBoomConfig.fir 383818:4]
  assign auto_client_out_a_bits_mask = inDes_io_out_bits_union; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 385:15 chipyard.TestHarness.SmallBoomConfig.fir 383821:4]
  assign auto_client_out_a_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 380:15 chipyard.TestHarness.SmallBoomConfig.fir 383819:4]
  assign auto_client_out_a_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 374:17 chipyard.TestHarness.SmallBoomConfig.fir 383813:4 Serdes.scala 382:17 chipyard.TestHarness.SmallBoomConfig.fir 383820:4]
  assign auto_client_out_d_ready = outArb_io_in_1_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383592:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383788:4]
  assign io_ser_in_ready = inDes_io_in_ready; // @[Serdes.scala 630:17 chipyard.TestHarness.SmallBoomConfig.fir 383809:4]
  assign io_ser_out_valid = outSer_io_out_valid; // @[Serdes.scala 627:16 chipyard.TestHarness.SmallBoomConfig.fir 383802:4]
  assign io_ser_out_bits = outSer_io_out_bits; // @[Serdes.scala 627:16 chipyard.TestHarness.SmallBoomConfig.fir 383801:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383515:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383516:4]
  assign monitor_io_in_a_ready = outArb_io_in_4_ready; // @[Serdes.scala 357:22 chipyard.TestHarness.SmallBoomConfig.fir 383735:4 Serdes.scala 625:18 chipyard.TestHarness.SmallBoomConfig.fir 383797:4]
  assign monitor_io_in_a_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_a_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_a_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_a_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_a_bits_source = auto_manager_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_a_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_a_bits_mask = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_a_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_d_ready = auto_manager_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign monitor_io_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 637:46 chipyard.TestHarness.SmallBoomConfig.fir 383877:4]
  assign monitor_io_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 461:15 chipyard.TestHarness.SmallBoomConfig.fir 383880:4]
  assign monitor_io_in_d_bits_param = inDes_io_out_bits_param[1:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 462:15 chipyard.TestHarness.SmallBoomConfig.fir 383881:4]
  assign monitor_io_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 463:15 chipyard.TestHarness.SmallBoomConfig.fir 383882:4]
  assign monitor_io_in_d_bits_source = inDes_io_out_bits_source[0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 464:15 chipyard.TestHarness.SmallBoomConfig.fir 383883:4]
  assign monitor_io_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[2:0]; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 468:17 chipyard.TestHarness.SmallBoomConfig.fir 383887:4]
  assign monitor_io_in_d_bits_denied = inDes_io_out_bits_union[0]; // @[Serdes.scala 469:30 chipyard.TestHarness.SmallBoomConfig.fir 383888:4]
  assign monitor_io_in_d_bits_corrupt = inDes_io_out_bits_corrupt; // @[Serdes.scala 460:17 chipyard.TestHarness.SmallBoomConfig.fir 383879:4 Serdes.scala 467:17 chipyard.TestHarness.SmallBoomConfig.fir 383885:4]
  assign outArb_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383546:4]
  assign outArb_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383547:4]
  assign outArb_io_in_1_valid = auto_client_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383510:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383537:4]
  assign outArb_io_in_1_bits_opcode = auto_client_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383510:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383537:4]
  assign outArb_io_in_1_bits_param = {{1'd0}, auto_client_out_d_bits_param}; // @[Serdes.scala 312:22 chipyard.TestHarness.SmallBoomConfig.fir 383594:4 Serdes.scala 315:20 chipyard.TestHarness.SmallBoomConfig.fir 383597:4]
  assign outArb_io_in_1_bits_size = {{1'd0}, auto_client_out_d_bits_size}; // @[Serdes.scala 312:22 chipyard.TestHarness.SmallBoomConfig.fir 383594:4 Serdes.scala 316:20 chipyard.TestHarness.SmallBoomConfig.fir 383598:4]
  assign outArb_io_in_1_bits_source = auto_client_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383510:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383537:4]
  assign outArb_io_in_1_bits_data = auto_client_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383510:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383537:4]
  assign outArb_io_in_1_bits_corrupt = auto_client_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 383510:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 383537:4]
  assign outArb_io_in_1_bits_union = {{6'd0}, _merged_bits_merged_union_T_1}; // @[Serdes.scala 312:22 chipyard.TestHarness.SmallBoomConfig.fir 383594:4 Serdes.scala 322:22 chipyard.TestHarness.SmallBoomConfig.fir 383604:4]
  assign outArb_io_in_1_bits_last = _merged_bits_last_last_T_2 | _merged_bits_last_last_T_3; // @[Edges.scala 231:37 chipyard.TestHarness.SmallBoomConfig.fir 383630:4]
  assign outArb_io_in_4_valid = auto_manager_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_opcode = auto_manager_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_param = auto_manager_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_size = auto_manager_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_source = {{3'd0}, auto_manager_in_a_bits_source}; // @[Serdes.scala 255:22 chipyard.TestHarness.SmallBoomConfig.fir 383737:4 Serdes.scala 260:20 chipyard.TestHarness.SmallBoomConfig.fir 383742:4]
  assign outArb_io_in_4_bits_address = auto_manager_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_data = auto_manager_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_corrupt = auto_manager_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_union = auto_manager_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 383512:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 383538:4]
  assign outArb_io_in_4_bits_last = _merged_bits_last_last_T_8 | _merged_bits_last_last_T_9; // @[Edges.scala 231:37 chipyard.TestHarness.SmallBoomConfig.fir 383773:4]
  assign outArb_io_out_ready = outSer_io_in_ready; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383800:4]
  assign outSer_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383549:4]
  assign outSer_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383550:4]
  assign outSer_io_in_valid = outArb_io_out_valid; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383799:4]
  assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_param = outArb_io_out_bits_param; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_size = outArb_io_out_bits_size; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_source = outArb_io_out_bits_source; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_address = outArb_io_out_bits_address; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_data = outArb_io_out_bits_data; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_corrupt = outArb_io_out_bits_corrupt; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_union = outArb_io_out_bits_union; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_in_bits_last = outArb_io_out_bits_last; // @[Serdes.scala 626:18 chipyard.TestHarness.SmallBoomConfig.fir 383798:4]
  assign outSer_io_out_ready = io_ser_out_ready; // @[Serdes.scala 627:16 chipyard.TestHarness.SmallBoomConfig.fir 383803:4]
  assign inDes_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 383805:4]
  assign inDes_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 383806:4]
  assign inDes_io_in_valid = io_ser_in_valid; // @[Serdes.scala 630:17 chipyard.TestHarness.SmallBoomConfig.fir 383808:4]
  assign inDes_io_in_bits = io_ser_in_bits; // @[Serdes.scala 630:17 chipyard.TestHarness.SmallBoomConfig.fir 383807:4]
  assign inDes_io_out_ready = _inDes_io_out_ready_T_8 ? 1'h0 : _inDes_io_out_ready_T_7; // @[Mux.scala 80:57 chipyard.TestHarness.SmallBoomConfig.fir 383924:4]
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383624:4]
      merged_bits_last_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383624:4]
    end else if (_merged_bits_last_T_1) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 383634:4]
      if (merged_bits_last_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 383635:6]
        if (merged_bits_last_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383623:4]
          merged_bits_last_counter_1 <= merged_bits_last_beats1_decode;
        end else begin
          merged_bits_last_counter_1 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_1 <= merged_bits_last_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383767:4]
      merged_bits_last_counter_4 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 383767:4]
    end else if (_merged_bits_last_T_4) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 383777:4]
      if (merged_bits_last_first_4) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 383778:6]
        if (merged_bits_last_beats1_opdata_3) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 383766:4]
          merged_bits_last_counter_4 <= merged_bits_last_beats1_decode_3;
        end else begin
          merged_bits_last_counter_4 <= 3'h0;
        end
      end else begin
        merged_bits_last_counter_4 <= merged_bits_last_counter1_4;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  merged_bits_last_counter_1 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  merged_bits_last_counter_4 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_54_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 383943:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 383944:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 383945:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
  input  [7:0]  io_in_d_bits_source // @[chipyard.TestHarness.SmallBoomConfig.fir 383946:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [639:0] _RAND_11;
  reg [639:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [639:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385437:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385744:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 383963:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 383969:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 383971:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 383972:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 383972:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 383973:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.SmallBoomConfig.fir 383974:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 383975:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 383976:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 383978:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 383979:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 383980:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 383981:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 383982:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 383984:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 383985:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 383987:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 383988:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 383989:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 383990:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 383991:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 383992:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 383993:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 383994:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 383995:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 383996:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 383997:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 383998:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 383999:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384000:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384001:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384002:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384003:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 384004:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 384005:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 384006:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384007:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384008:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384009:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384010:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384011:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384012:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384013:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384014:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384015:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384016:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384017:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384018:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384019:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384020:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384021:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384022:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384023:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384024:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384025:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384026:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384027:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 384028:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 384029:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 384030:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 384037:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 384060:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 384076:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 384077:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 384079:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 384080:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384086:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384111:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384112:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384119:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384120:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384126:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384127:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 384132:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384134:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384135:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 384140:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 384141:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384143:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384144:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 384149:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384151:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384152:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 384158:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 384238:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384240:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384241:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 384264:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384298:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384299:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 384318:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384320:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384321:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 384326:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384328:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384329:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 384343:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 384369:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384371:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384372:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 384408:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 384464:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 384465:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 384466:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384468:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384469:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 384475:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 384520:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384522:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384523:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 384537:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 384582:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384584:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384585:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 384599:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 384644:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384646:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384647:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 384671:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384673:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384674:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 384685:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 384691:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384694:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384695:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 384700:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384702:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384703:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 384733:6]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 384791:6]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 384850:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 384885:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 384921:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 384987:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 384996:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 384998:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 384999:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 385010:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 385011:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 385012:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 385013:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 385014:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 385015:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 385016:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 385018:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385020:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385021:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 385026:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385028:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385029:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 385034:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385036:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385037:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 385042:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385044:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385045:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 385050:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385052:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385053:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 385060:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 385068:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385076:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385078:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385079:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 385090:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 385092:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 385093:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 385096:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 385097:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 385099:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385101:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385102:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 385115:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385117:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385118:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 385123:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385125:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385126:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 385149:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 385158:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 385159:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 385160:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385170:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385172:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385173:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385192:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385194:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385195:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 385216:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 385216:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 385217:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 385221:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 385222:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 385222:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 385223:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 385228:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 385233:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 385234:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 385258:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 385261:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 385260:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 385262:6 chipyard.TestHarness.SmallBoomConfig.fir 385209:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 385265:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 385270:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 385271:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 385273:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 385274:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 385276:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 385276:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385267:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 385272:6 chipyard.TestHarness.SmallBoomConfig.fir 385255:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 385277:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 385277:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385267:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 385275:6 chipyard.TestHarness.SmallBoomConfig.fir 385257:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 385280:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 385280:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 385282:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 385284:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385286:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385287:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385267:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 385269:6 chipyard.TestHarness.SmallBoomConfig.fir 385207:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385267:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 385278:6 chipyard.TestHarness.SmallBoomConfig.fir 385211:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 385267:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 385281:6 chipyard.TestHarness.SmallBoomConfig.fir 385213:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 385302:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 385304:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 385305:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 385307:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 385306:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 385308:6 chipyard.TestHarness.SmallBoomConfig.fir 385296:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 385311:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 385314:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 385323:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 385323:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 385315:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 385317:6 chipyard.TestHarness.SmallBoomConfig.fir 385294:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 385315:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 385324:6 chipyard.TestHarness.SmallBoomConfig.fir 385298:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 385340:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 385341:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 385342:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 385344:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385346:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385347:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 385353:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385354:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385354:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385354:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385354:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 385354:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 385355:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385357:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385358:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 385363:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385365:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385366:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385214:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 385224:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 385374:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385376:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385376:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385376:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385376:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 385376:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 385377:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385379:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385380:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385225:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 385235:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 385385:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 385385:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385387:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385388:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 385396:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 385397:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 385399:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 385401:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 385403:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 385404:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385406:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385407:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385208:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385295:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 385413:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 385414:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 385415:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 385416:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385418:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385419:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385206:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 385424:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385293:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 385425:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 385426:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385210:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 385428:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385297:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 385429:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 385430:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385212:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 385432:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 385434:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 385436:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 385439:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 385440:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 385441:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 385442:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 385443:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 385444:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385446:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385447:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 385453:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 385457:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 385461:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 385463:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385498:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 385500:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 385501:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 385534:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 385539:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 385540:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 385618:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 385620:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 385626:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 385628:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 385629:4 Monitor.scala 784:21 chipyard.TestHarness.SmallBoomConfig.fir 385631:6 chipyard.TestHarness.SmallBoomConfig.fir 385610:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 385629:4 Monitor.scala 785:21 chipyard.TestHarness.SmallBoomConfig.fir 385638:6 chipyard.TestHarness.SmallBoomConfig.fir 385614:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 385664:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385668:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385669:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385522:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 385541:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 385687:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385689:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385690:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385609:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.SmallBoomConfig.fir 385732:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.SmallBoomConfig.fir 385733:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 385613:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.SmallBoomConfig.fir 385736:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 385741:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 385743:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.SmallBoomConfig.fir 385746:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.SmallBoomConfig.fir 385747:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.SmallBoomConfig.fir 385748:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.SmallBoomConfig.fir 385749:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.SmallBoomConfig.fir 385750:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.SmallBoomConfig.fir 385751:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385753:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385754:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.SmallBoomConfig.fir 385760:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384088:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384186:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384283:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384374:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384439:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384503:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384565:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384627:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384697:10]
  wire  _GEN_202 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384739:10]
  wire  _GEN_208 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384797:10]
  wire  _GEN_214 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384856:10]
  wire  _GEN_216 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384891:10]
  wire  _GEN_218 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384927:10]
  wire  _GEN_220 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385360:10]
  wire  _GEN_225 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385382:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385437:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 385744:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 384996:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 384996:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385006:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385007:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385061:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 385062:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385061:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 385063:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385061:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 385064:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385061:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 385065:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 385061:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 385066:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385076:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385076:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385086:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385087:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 385150:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 385151:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 385150:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 385153:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 385150:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 385154:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 385158:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 385158:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 385427:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 385159:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 385159:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 385431:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 385160:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 385160:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 385435:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385170:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385170:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385180:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385181:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385192:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385192:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385202:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385203:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 385436:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 385436:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 385458:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 385459:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 385454:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 385461:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 385461:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.SmallBoomConfig.fir 385734:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 385463:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 385463:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 385742:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385498:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 385498:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 385508:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 385509:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 385743:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 385743:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.SmallBoomConfig.fir 385767:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.SmallBoomConfig.fir 385768:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.SmallBoomConfig.fir 385761:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384088:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384089:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384107:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384108:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384114:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384115:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384122:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384123:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384129:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384130:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384137:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384138:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384146:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384147:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384154:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384155:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384186:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384187:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384205:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384206:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384212:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384213:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384220:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384221:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384227:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384228:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384235:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384236:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384243:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384244:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384252:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384253:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384260:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384261:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384283:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384284:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384301:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384302:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384308:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384309:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384315:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384316:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384323:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384324:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384331:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384332:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384339:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384340:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384374:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384375:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384381:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384382:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384388:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384389:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384396:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384397:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384404:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384405:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384439:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384440:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384446:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384447:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384453:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384454:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384461:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384462:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384471:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384472:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384503:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384504:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384510:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384511:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384517:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384518:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384525:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384526:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384533:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384534:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384565:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384566:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384572:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384573:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384579:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384580:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384587:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384588:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384595:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384596:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384627:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384628:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384634:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384635:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384641:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384642:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384649:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384650:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384657:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384658:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384665:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 384666:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384676:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384677:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384697:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384698:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384705:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384706:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384739:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384740:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384746:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384747:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384754:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_202 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384755:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384797:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384798:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384804:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384805:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384812:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384813:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384856:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_214 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384857:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384891:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_216 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384892:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384927:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_218 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 384928:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385023:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385024:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385031:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385032:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385039:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385040:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385047:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385048:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385055:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385056:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385104:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385105:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385120:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385121:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385128:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385129:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385289:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385290:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385349:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385350:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385360:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385361:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385368:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_220 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385369:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385382:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385383:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385390:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_225 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385391:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385409:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385410:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385421:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385422:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385449:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385450:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385671:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385672:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385692:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 385693:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:31)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385756:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 385757:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  size_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  source_1 = _RAND_9[7:0];
  _RAND_10 = {5{`RANDOM}};
  inflight = _RAND_10[159:0];
  _RAND_11 = {20{`RANDOM}};
  inflight_opcodes = _RAND_11[639:0];
  _RAND_12 = {20{`RANDOM}};
  inflight_sizes = _RAND_12[639:0];
  _RAND_13 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  watchdog = _RAND_15[31:0];
  _RAND_16 = {5{`RANDOM}};
  inflight_1 = _RAND_16[159:0];
  _RAND_17 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_17[639:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  watchdog_1 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLRAM_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 385771:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 385772:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 385773:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input  [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  output [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
  output [63:0] auto_in_d_bits_data // @[chipyard.TestHarness.SmallBoomConfig.fir 385774:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
  wire [8:0] mem_RW0_addr; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_en; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_clk; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmode; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_wdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire [7:0] mem_RW0_rdata_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_0; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_1; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_2; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_3; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_4; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_5; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_6; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  wire  mem_RW0_wmask_7; // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
  reg  r_full; // @[SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385820:4]
  reg [1:0] r_size; // @[SRAM.scala 137:26 chipyard.TestHarness.SmallBoomConfig.fir 385823:4]
  reg [7:0] r_source; // @[SRAM.scala 138:26 chipyard.TestHarness.SmallBoomConfig.fir 385824:4]
  reg  r_read; // @[SRAM.scala 139:26 chipyard.TestHarness.SmallBoomConfig.fir 385825:4]
  reg  REG; // @[SRAM.scala 321:58 chipyard.TestHarness.SmallBoomConfig.fir 386345:4]
  reg [7:0] r_1; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_1 = REG ? mem_RW0_rdata_1 : r_1; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  reg [7:0] r_0; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_0 = REG ? mem_RW0_rdata_0 : r_0; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  reg [7:0] r_3; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_3 = REG ? mem_RW0_rdata_3 : r_3; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  reg [7:0] r_2; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_2 = REG ? mem_RW0_rdata_2 : r_2; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  wire [31:0] r_corrected_lo = {r_raw_data_3,r_raw_data_2,r_raw_data_1,r_raw_data_0}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 385888:4]
  reg [7:0] r_5; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_5 = REG ? mem_RW0_rdata_5 : r_5; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  reg [7:0] r_4; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_4 = REG ? mem_RW0_rdata_4 : r_4; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  reg [7:0] r_7; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_7 = REG ? mem_RW0_rdata_7 : r_7; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  reg [7:0] r_6; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 386347:4]
  wire [7:0] r_raw_data_6 = REG ? mem_RW0_rdata_6 : r_6; // @[package.scala 79:42 chipyard.TestHarness.SmallBoomConfig.fir 386358:4]
  wire [31:0] r_corrected_hi = {r_raw_data_7,r_raw_data_6,r_raw_data_5,r_raw_data_4}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 385891:4]
  wire  _bundleIn_0_a_ready_T_2 = ~r_full; // @[SRAM.scala 243:41 chipyard.TestHarness.SmallBoomConfig.fir 386071:4]
  wire  in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.SmallBoomConfig.fir 386072:4]
  wire  a_read = auto_in_a_bits_opcode == 3'h4; // @[SRAM.scala 251:35 chipyard.TestHarness.SmallBoomConfig.fir 386080:4]
  wire  _GEN_22 = auto_in_d_ready ? 1'h0 : r_full; // @[SRAM.scala 273:20 chipyard.TestHarness.SmallBoomConfig.fir 386109:4 SRAM.scala 273:29 chipyard.TestHarness.SmallBoomConfig.fir 386110:6 SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385820:4]
  wire  _T_18 = in_a_ready & auto_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 386112:4]
  wire  _T_19 = ~a_read; // @[SRAM.scala 287:13 chipyard.TestHarness.SmallBoomConfig.fir 386126:6]
  wire  _GEN_24 = _T_18 | _GEN_22; // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386113:4 SRAM.scala 275:18 chipyard.TestHarness.SmallBoomConfig.fir 386114:6]
  wire  a_lanes_lo_lo_lo = |auto_in_a_bits_mask[0]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386250:4]
  wire  a_lanes_lo_lo_hi = |auto_in_a_bits_mask[1]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386252:4]
  wire  a_lanes_lo_hi_lo = |auto_in_a_bits_mask[2]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386254:4]
  wire  a_lanes_lo_hi_hi = |auto_in_a_bits_mask[3]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386256:4]
  wire  a_lanes_hi_lo_lo = |auto_in_a_bits_mask[4]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386258:4]
  wire  a_lanes_hi_lo_hi = |auto_in_a_bits_mask[5]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386260:4]
  wire  a_lanes_hi_hi_lo = |auto_in_a_bits_mask[6]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386262:4]
  wire  a_lanes_hi_hi_hi = |auto_in_a_bits_mask[7]; // @[SRAM.scala 303:95 chipyard.TestHarness.SmallBoomConfig.fir 386264:4]
  wire [7:0] a_lanes = {a_lanes_hi_hi_hi,a_lanes_hi_hi_lo,a_lanes_hi_lo_hi,a_lanes_hi_lo_lo,a_lanes_lo_hi_hi,
    a_lanes_lo_hi_lo,a_lanes_lo_lo_hi,a_lanes_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386271:4]
  wire  wen = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.SmallBoomConfig.fir 386279:4]
  wire  _ren_T = ~wen; // @[SRAM.scala 310:15 chipyard.TestHarness.SmallBoomConfig.fir 386282:4]
  wire  ren = _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.SmallBoomConfig.fir 386284:4]
  wire  index_lo_lo_lo = auto_in_a_bits_address[3]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386303:4]
  wire  index_lo_lo_hi = auto_in_a_bits_address[4]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386304:4]
  wire  index_lo_hi_lo = auto_in_a_bits_address[5]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386305:4]
  wire  index_lo_hi_hi = auto_in_a_bits_address[6]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386306:4]
  wire  index_hi_lo_lo = auto_in_a_bits_address[7]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386307:4]
  wire  index_hi_lo_hi = auto_in_a_bits_address[8]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386308:4]
  wire  index_hi_hi_lo = auto_in_a_bits_address[9]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386309:4]
  wire  index_hi_hi_hi_lo = auto_in_a_bits_address[10]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386310:4]
  wire  index_hi_hi_hi_hi = auto_in_a_bits_address[11]; // @[SRAM.scala 320:60 chipyard.TestHarness.SmallBoomConfig.fir 386311:4]
  wire [3:0] index_lo = {index_lo_hi_hi,index_lo_hi_lo,index_lo_lo_hi,index_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386331:4]
  wire [4:0] index_hi = {index_hi_hi_hi_hi,index_hi_hi_hi_lo,index_hi_hi_lo,index_hi_lo_hi,index_hi_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386335:4]
  TLMonitor_54_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 385781:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source)
  );



  mem_inTestHarness mem ( // @[DescribedSRAM.scala 19:26 chipyard.TestHarness.SmallBoomConfig.fir 385805:4]
    .RW0_addr(mem_RW0_addr),
    .RW0_en(mem_RW0_en),
    .RW0_clk(mem_RW0_clk),
    .RW0_wmode(mem_RW0_wmode),
    .RW0_wdata_0(mem_RW0_wdata_0),
    .RW0_wdata_1(mem_RW0_wdata_1),
    .RW0_wdata_2(mem_RW0_wdata_2),
    .RW0_wdata_3(mem_RW0_wdata_3),
    .RW0_wdata_4(mem_RW0_wdata_4),
    .RW0_wdata_5(mem_RW0_wdata_5),
    .RW0_wdata_6(mem_RW0_wdata_6),
    .RW0_wdata_7(mem_RW0_wdata_7),
    .RW0_rdata_0(mem_RW0_rdata_0),
    .RW0_rdata_1(mem_RW0_rdata_1),
    .RW0_rdata_2(mem_RW0_rdata_2),
    .RW0_rdata_3(mem_RW0_rdata_3),
    .RW0_rdata_4(mem_RW0_rdata_4),
    .RW0_rdata_5(mem_RW0_rdata_5),
    .RW0_rdata_6(mem_RW0_rdata_6),
    .RW0_rdata_7(mem_RW0_rdata_7),
    .RW0_wmask_0(mem_RW0_wmask_0),
    .RW0_wmask_1(mem_RW0_wmask_1),
    .RW0_wmask_2(mem_RW0_wmask_2),
    .RW0_wmask_3(mem_RW0_wmask_3),
    .RW0_wmask_4(mem_RW0_wmask_4),
    .RW0_wmask_5(mem_RW0_wmask_5),
    .RW0_wmask_6(mem_RW0_wmask_6),
    .RW0_wmask_7(mem_RW0_wmask_7)
  );
  assign auto_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.SmallBoomConfig.fir 386072:4]
  assign auto_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.SmallBoomConfig.fir 386051:4]
  assign auto_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 SRAM.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 385999:4]
  assign auto_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.SmallBoomConfig.fir 386001:4]
  assign auto_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.SmallBoomConfig.fir 386003:4]
  assign auto_in_d_bits_data = {r_corrected_hi,r_corrected_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 385899:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 385782:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 385783:4]
  assign monitor_io_in_a_ready = _bundleIn_0_a_ready_T_2 | auto_in_d_ready; // @[SRAM.scala 243:49 chipyard.TestHarness.SmallBoomConfig.fir 386072:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 385804:4]
  assign monitor_io_in_d_valid = r_full; // @[SRAM.scala 240:65 chipyard.TestHarness.SmallBoomConfig.fir 386051:4]
  assign monitor_io_in_d_bits_opcode = {{2'd0}, r_read}; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 385779:4 SRAM.scala 209:23 chipyard.TestHarness.SmallBoomConfig.fir 385999:4]
  assign monitor_io_in_d_bits_size = r_size; // @[SRAM.scala 211:29 chipyard.TestHarness.SmallBoomConfig.fir 386001:4]
  assign monitor_io_in_d_bits_source = r_source; // @[SRAM.scala 212:29 chipyard.TestHarness.SmallBoomConfig.fir 386003:4]
  assign mem_RW0_wdata_0 = auto_in_a_bits_data[7:0]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386131:4]
  assign mem_RW0_wdata_1 = auto_in_a_bits_data[15:8]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386132:4]
  assign mem_RW0_wdata_2 = auto_in_a_bits_data[23:16]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386133:4]
  assign mem_RW0_wdata_3 = auto_in_a_bits_data[31:24]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386134:4]
  assign mem_RW0_wdata_4 = auto_in_a_bits_data[39:32]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386135:4]
  assign mem_RW0_wdata_5 = auto_in_a_bits_data[47:40]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386136:4]
  assign mem_RW0_wdata_6 = auto_in_a_bits_data[55:48]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386137:4]
  assign mem_RW0_wdata_7 = auto_in_a_bits_data[63:56]; // @[SRAM.scala 291:67 chipyard.TestHarness.SmallBoomConfig.fir 386138:4]
  assign mem_RW0_wmask_0 = a_lanes[0]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386368:6]
  assign mem_RW0_wmask_1 = a_lanes[1]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386369:6]
  assign mem_RW0_wmask_2 = a_lanes[2]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386370:6]
  assign mem_RW0_wmask_3 = a_lanes[3]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386371:6]
  assign mem_RW0_wmask_4 = a_lanes[4]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386372:6]
  assign mem_RW0_wmask_5 = a_lanes[5]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386373:6]
  assign mem_RW0_wmask_6 = a_lanes[6]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386374:6]
  assign mem_RW0_wmask_7 = a_lanes[7]; // @[SRAM.scala 322:46 chipyard.TestHarness.SmallBoomConfig.fir 386375:6]
  assign mem_RW0_wmode = _T_18 & _T_19; // @[SRAM.scala 309:52 chipyard.TestHarness.SmallBoomConfig.fir 386279:4]
  assign mem_RW0_clk = clock;
  assign mem_RW0_en = ren | wen;
  assign mem_RW0_addr = {index_hi,index_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 386336:4]
  always @(posedge clock) begin
    if (reset) begin // @[SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385820:4]
      r_full <= 1'h0; // @[SRAM.scala 134:30 chipyard.TestHarness.SmallBoomConfig.fir 385820:4]
    end else begin
      r_full <= _GEN_24;
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386113:4]
      r_size <= auto_in_a_bits_size; // @[SRAM.scala 279:18 chipyard.TestHarness.SmallBoomConfig.fir 386118:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386113:4]
      r_source <= auto_in_a_bits_source; // @[SRAM.scala 280:18 chipyard.TestHarness.SmallBoomConfig.fir 386119:6]
    end
    if (_T_18) begin // @[SRAM.scala 274:24 chipyard.TestHarness.SmallBoomConfig.fir 386113:4]
      r_read <= a_read; // @[SRAM.scala 281:18 chipyard.TestHarness.SmallBoomConfig.fir 386120:6]
    end
    REG <= _ren_T & _T_18; // @[SRAM.scala 310:20 chipyard.TestHarness.SmallBoomConfig.fir 386284:4]
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_1 <= mem_RW0_rdata_1; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386350:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_0 <= mem_RW0_rdata_0; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386349:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_3 <= mem_RW0_rdata_3; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386352:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_2 <= mem_RW0_rdata_2; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386351:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_5 <= mem_RW0_rdata_5; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386354:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_4 <= mem_RW0_rdata_4; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386353:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_7 <= mem_RW0_rdata_7; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386356:6]
    end
    if (REG) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 386348:4]
      r_6 <= mem_RW0_rdata_6; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 386355:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_size = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r_source = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  r_read = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r_5 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  r_4 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  r_7 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_6 = _RAND_12[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar_10_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 386412:2]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [2:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [3:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [2:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [3:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 386415:4]
);
  assign auto_in_a_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386420:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386424:4]
  assign auto_in_d_valid = auto_out_d_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.SmallBoomConfig.fir 386836:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386420:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386424:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386420:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386424:4]
  assign auto_in_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386420:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386424:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source; // @[Xbar.scala 228:69 chipyard.TestHarness.SmallBoomConfig.fir 386535:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Xbar.scala 323:53 chipyard.TestHarness.SmallBoomConfig.fir 386597:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386420:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386424:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386420:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386424:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 386420:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 386424:4]
  assign auto_out_a_valid = auto_in_a_valid; // @[ReadyValidCancel.scala 21:38 chipyard.TestHarness.SmallBoomConfig.fir 386861:4]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
  assign auto_out_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Xbar.scala 237:55 chipyard.TestHarness.SmallBoomConfig.fir 386489:4]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
  assign auto_out_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
  assign auto_out_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
  assign auto_out_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 386422:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 386425:4]
endmodule
module TLMonitor_55_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 386938:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 386939:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 386940:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [1:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [7:0]  io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [1:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input  [7:0]  io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 386941:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [639:0] _RAND_14;
  reg [639:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [639:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388432:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388739:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 386958:6]
  wire [5:0] _is_aligned_mask_T_1 = 6'h7 << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 386964:6]
  wire [2:0] is_aligned_mask = ~_is_aligned_mask_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 386966:6]
  wire [28:0] _GEN_71 = {{26'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 386967:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 386967:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 386968:6]
  wire [2:0] _mask_sizeOH_T = {{1'd0}, io_in_a_bits_size}; // @[Misc.scala 201:34 chipyard.TestHarness.SmallBoomConfig.fir 386969:6]
  wire [1:0] mask_sizeOH_shiftAmount = _mask_sizeOH_T[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 386970:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 386971:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 386973:6]
  wire  _mask_T = io_in_a_bits_size >= 2'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 386974:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 386975:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 386976:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 386977:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 386979:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 386980:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 386982:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 386983:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 386984:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 386985:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 386986:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 386987:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 386988:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 386989:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 386990:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 386991:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 386992:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 386993:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 386994:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 386995:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 386996:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 386997:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 386998:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 386999:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 387000:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 387001:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387002:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387003:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387004:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387005:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387006:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387007:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387008:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387009:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387010:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387011:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387012:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387013:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387014:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387015:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387016:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387017:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387018:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387019:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387020:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387021:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387022:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 387023:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 387024:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 387025:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 387032:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 387055:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 387071:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 387072:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 387074:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 387075:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387081:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387106:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387107:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387114:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387115:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387121:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387122:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 387127:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387129:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387130:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 387135:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 387136:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387138:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387139:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 387144:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387146:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387147:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 387153:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 387233:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387235:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387236:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 387259:6]
  wire  _T_175 = _T_37 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387293:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387294:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 387313:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387315:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387316:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 387321:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387323:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387324:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 387338:6]
  wire  _T_218 = _source_ok_T_4 & _T_37; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 387364:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387366:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387367:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 387403:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 387459:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 387460:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 387461:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387463:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387464:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 387470:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 387515:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387517:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387518:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 387532:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 387577:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387579:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387580:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 387594:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 387639:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387641:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387642:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 387666:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387668:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387669:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 8'h9f; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 387680:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 387686:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387689:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387690:8]
  wire  _T_405 = io_in_d_bits_size >= 2'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 387695:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387697:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387698:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 387703:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387705:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387706:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 387711:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387713:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387714:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 387719:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387721:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387722:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 387728:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 387752:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387754:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387755:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 387760:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387762:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387763:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 387786:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 387827:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387829:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387830:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 387845:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 387880:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 387916:6]
  wire  a_first_done = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 387982:4]
  reg  a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 387991:4]
  wire  a_first_counter1 = a_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 387993:4]
  wire  a_first = ~a_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 387994:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 388005:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 388006:4]
  reg [1:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 388007:4]
  reg [7:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 388008:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 388009:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 388010:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 388011:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 388013:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388015:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388016:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 388021:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388023:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388024:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 388029:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388031:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388032:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 388037:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388039:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388040:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 388045:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388047:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388048:6]
  wire  _T_565 = a_first_done & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 388055:4]
  wire  d_first_done = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 388063:4]
  reg  d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388071:4]
  wire  d_first_counter1 = d_first_counter - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388073:4]
  wire  d_first = ~d_first_counter; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388074:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 388085:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 388086:4]
  reg [1:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 388087:4]
  reg [7:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 388088:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 388089:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 388090:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 388091:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 388092:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 388094:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388096:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388097:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 388102:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388104:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388105:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 388110:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388112:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388113:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 388118:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388120:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388121:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 388126:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388128:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388129:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 388134:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388136:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388137:6]
  wire  _T_593 = d_first_done & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 388144:4]
  reg [159:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 388153:4]
  reg [639:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 388154:4]
  reg [639:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 388155:4]
  reg  a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388165:4]
  wire  a_first_counter1_1 = a_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388167:4]
  wire  a_first_1 = ~a_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388168:4]
  reg  d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388187:4]
  wire  d_first_counter1_1 = d_first_counter_1 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388189:4]
  wire  d_first_1 = ~d_first_counter_1; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388190:4]
  wire [9:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 388211:4]
  wire [10:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 388211:4]
  wire [639:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 388212:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 388216:4]
  wire [639:0] _GEN_73 = {{624'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 388217:4]
  wire [639:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 388217:4]
  wire [639:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[639:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 388218:4]
  wire [639:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 388223:4]
  wire [639:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 388228:4]
  wire [639:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[639:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 388229:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 388253:4]
  wire [255:0] _a_set_wo_ready_T = 256'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 388256:6]
  wire [255:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 388255:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 388257:6 chipyard.TestHarness.SmallBoomConfig.fir 388204:4]
  wire  _T_597 = a_first_done & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 388260:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 388265:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 388266:6]
  wire [2:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 388268:6]
  wire [2:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 3'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 388269:6]
  wire [9:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 388271:6]
  wire [10:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 388271:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388262:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 388267:6 chipyard.TestHarness.SmallBoomConfig.fir 388250:4]
  wire [2050:0] _GEN_79 = {{2047'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 388272:6]
  wire [2050:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 388272:6]
  wire [2:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 3'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388262:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 388270:6 chipyard.TestHarness.SmallBoomConfig.fir 388252:4]
  wire [2049:0] _GEN_81 = {{2047'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 388275:6]
  wire [2049:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 388275:6]
  wire [159:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 388277:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 388279:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388281:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388282:6]
  wire [255:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 256'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388262:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 388264:6 chipyard.TestHarness.SmallBoomConfig.fir 388202:4]
  wire [2050:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 2051'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388262:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 388273:6 chipyard.TestHarness.SmallBoomConfig.fir 388206:4]
  wire [2049:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 2050'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 388262:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 388276:6 chipyard.TestHarness.SmallBoomConfig.fir 388208:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 388297:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 388299:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 388300:4]
  wire [255:0] _d_clr_wo_ready_T = 256'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 388302:6]
  wire [255:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 388301:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 388303:6 chipyard.TestHarness.SmallBoomConfig.fir 388291:4]
  wire  _T_610 = d_first_done & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 388306:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 388309:4]
  wire [2062:0] _GEN_83 = {{2047'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 388318:6]
  wire [2062:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 388318:6]
  wire [255:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 388310:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 388312:6 chipyard.TestHarness.SmallBoomConfig.fir 388289:4]
  wire [2062:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 388310:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 388319:6 chipyard.TestHarness.SmallBoomConfig.fir 388293:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 388335:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 388336:6]
  wire [159:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 388337:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 388339:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388341:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388342:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 388348:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388349:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388349:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388349:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388349:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 388349:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 388350:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388352:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388353:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 388358:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388360:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388361:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388209:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 388219:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 388369:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388371:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388371:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388371:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388371:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 388371:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 388372:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388374:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388375:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388220:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 388230:4]
  wire [3:0] _GEN_86 = {{2'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 388380:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 388380:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388382:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388383:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 388391:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 388392:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 388394:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 388396:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 388398:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 388399:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388401:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388402:6]
  wire [159:0] a_set_wo_ready = _GEN_15[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388203:4]
  wire [159:0] d_clr_wo_ready = _GEN_21[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388290:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 388408:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 388409:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 388410:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 388411:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388413:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388414:4]
  wire [159:0] a_set = _GEN_16[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388201:4]
  wire [159:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 388419:4]
  wire [159:0] d_clr = _GEN_22[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388288:4]
  wire [159:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 388420:4]
  wire [159:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 388421:4]
  wire [639:0] a_opcodes_set = _GEN_19[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388205:4]
  wire [639:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 388423:4]
  wire [639:0] d_opcodes_clr = _GEN_23[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388292:4]
  wire [639:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 388424:4]
  wire [639:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 388425:4]
  wire [639:0] a_sizes_set = _GEN_20[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388207:4]
  wire [639:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 388427:4]
  wire [639:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 388429:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 388431:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 388434:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 388435:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 388436:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 388437:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 388438:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 388439:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388441:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388442:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 388448:4]
  wire  _T_676 = a_first_done | d_first_done; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 388452:4]
  reg [159:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 388456:4]
  reg [639:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 388458:4]
  reg  d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388493:4]
  wire  d_first_counter1_2 = d_first_counter_2 - 1'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 388495:4]
  wire  d_first_2 = ~d_first_counter_2; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 388496:4]
  wire [639:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 388529:4]
  wire [639:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 388534:4]
  wire [639:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[639:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 388535:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 388613:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 388615:4]
  wire  _T_698 = d_first_done & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 388621:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 388623:4]
  wire [255:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 256'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 388624:4 Monitor.scala 784:21 chipyard.TestHarness.SmallBoomConfig.fir 388626:6 chipyard.TestHarness.SmallBoomConfig.fir 388605:4]
  wire [2062:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 2063'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 388624:4 Monitor.scala 785:21 chipyard.TestHarness.SmallBoomConfig.fir 388633:6 chipyard.TestHarness.SmallBoomConfig.fir 388609:4]
  wire [159:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 388659:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388663:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388664:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388517:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 388536:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 388682:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388684:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388685:8]
  wire [159:0] d_clr_1 = _GEN_67[159:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388604:4]
  wire [159:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.SmallBoomConfig.fir 388727:4]
  wire [159:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.SmallBoomConfig.fir 388728:4]
  wire [639:0] d_opcodes_clr_1 = _GEN_68[639:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 388608:4]
  wire [639:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.SmallBoomConfig.fir 388731:4]
  wire [639:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 388736:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 388738:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.SmallBoomConfig.fir 388741:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.SmallBoomConfig.fir 388742:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.SmallBoomConfig.fir 388743:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.SmallBoomConfig.fir 388744:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.SmallBoomConfig.fir 388745:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.SmallBoomConfig.fir 388746:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388748:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388749:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.SmallBoomConfig.fir 388755:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387083:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387181:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387278:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387369:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387434:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387498:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387560:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387622:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387692:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387734:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387792:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387851:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387886:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387922:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388355:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388377:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388432:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 388739:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 387991:4]
      a_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 387991:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388001:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388002:6]
        a_first_counter <= 1'h0;
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388056:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 388057:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388056:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 388058:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388056:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 388059:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388056:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 388060:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 388056:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 388061:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388071:4]
      d_first_counter <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388071:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388081:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388082:6]
        d_first_counter <= 1'h0;
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388145:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 388146:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388145:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 388147:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388145:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 388148:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388145:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 388149:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388145:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 388150:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 388145:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 388151:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 388153:4]
      inflight <= 160'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 388153:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 388422:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 388154:4]
      inflight_opcodes <= 640'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 388154:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 388426:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 388155:4]
      inflight_sizes <= 640'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 388155:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 388430:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388165:4]
      a_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388165:4]
    end else if (a_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388175:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388176:6]
        a_first_counter_1 <= 1'h0;
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388187:4]
      d_first_counter_1 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388187:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388197:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388198:6]
        d_first_counter_1 <= 1'h0;
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 388431:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 388431:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 388453:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 388454:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 388449:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 388456:4]
      inflight_1 <= 160'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 388456:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.SmallBoomConfig.fir 388729:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 388458:4]
      inflight_sizes_1 <= 640'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 388458:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 388737:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388493:4]
      d_first_counter_2 <= 1'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 388493:4]
    end else if (d_first_done) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 388503:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 388504:6]
        d_first_counter_2 <= 1'h0;
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 388738:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 388738:4]
    end else if (d_first_done) begin // @[Monitor.scala 819:47 chipyard.TestHarness.SmallBoomConfig.fir 388762:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.SmallBoomConfig.fir 388763:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.SmallBoomConfig.fir 388756:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387083:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387084:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387102:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387103:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387109:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387110:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387117:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387118:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387124:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387125:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387132:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387133:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387141:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387142:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387149:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387150:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387181:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387182:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387200:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387201:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387207:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387208:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387215:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387216:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387222:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387223:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387230:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387231:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387238:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387239:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387247:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387248:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387255:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387256:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387278:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387279:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387296:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387297:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387303:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387304:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387310:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387311:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387318:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387319:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387326:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387327:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387334:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387335:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387369:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387370:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387376:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387377:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387383:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387384:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387391:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387392:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387399:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387400:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387434:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387435:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387441:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387442:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387448:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387449:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387456:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387457:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387466:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387467:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387498:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387499:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387505:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387506:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387512:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387513:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387520:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387521:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387528:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387529:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387560:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387561:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387567:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387568:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387574:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387575:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387582:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387583:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387590:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387591:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387622:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387623:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387629:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387630:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387636:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387637:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387644:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387645:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387652:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387653:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387660:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 387661:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387671:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387672:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387692:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387693:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387700:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387701:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387708:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387709:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387716:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387717:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387724:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387725:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387734:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387735:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387741:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387742:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387749:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387750:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387757:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387758:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387765:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387766:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387773:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387774:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387782:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387783:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387792:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387793:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387799:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387800:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387807:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387808:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387815:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387816:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387823:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387824:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387832:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387833:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387841:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387842:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387851:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387852:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387859:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387860:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387867:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387868:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387876:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387877:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387886:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387887:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387894:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387895:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387903:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387904:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387912:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387913:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387922:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387923:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387930:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387931:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387938:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387939:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387947:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 387948:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388018:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388019:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388026:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388027:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388034:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388035:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388042:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388043:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388050:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388051:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388099:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388100:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388107:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388108:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388115:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388116:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388123:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388124:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388131:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388132:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388139:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388140:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388284:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388285:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388344:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388345:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388355:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388356:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388363:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388364:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388377:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388378:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388385:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388386:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388404:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388405:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388416:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388417:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388444:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388445:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388666:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388667:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388687:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 388688:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:45)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388751:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 388752:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {5{`RANDOM}};
  inflight = _RAND_13[159:0];
  _RAND_14 = {20{`RANDOM}};
  inflight_opcodes = _RAND_14[639:0];
  _RAND_15 = {20{`RANDOM}};
  inflight_sizes = _RAND_15[639:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {5{`RANDOM}};
  inflight_1 = _RAND_19[159:0];
  _RAND_20 = {20{`RANDOM}};
  inflight_sizes_1 = _RAND_20[639:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_44_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 388766:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 388767:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 388768:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input  [1:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input  [7:0]  io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input  [63:0] io_enq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output [1:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output [7:0]  io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output [63:0] io_deq_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 388769:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_opcode [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [2:0] ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_opcode_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [2:0] ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_opcode_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_opcode_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_opcode_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg [2:0] ram_param [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [2:0] ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_param_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [2:0] ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_param_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_param_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_param_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg [1:0] ram_size [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [1:0] ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_size_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [1:0] ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_size_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_size_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_size_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg [7:0] ram_source [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [7:0] ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_source_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [7:0] ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_source_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_source_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_source_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg [28:0] ram_address [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [28:0] ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_address_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [28:0] ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_address_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_address_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_address_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg [7:0] ram_mask [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [7:0] ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_mask_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [7:0] ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_mask_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_mask_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_mask_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg [63:0] ram_data [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [63:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire [63:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_data_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg  ram_corrupt [0:1]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_corrupt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_corrupt_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_corrupt_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  wire  ram_corrupt_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  reg  value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388772:4]
  reg  value_1; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388773:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 388774:4]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 388775:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 388776:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 388777:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 388778:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 388779:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 388782:4]
  wire  _value_T_1 = value + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 388797:6]
  wire  _value_T_3 = value_1 + 1'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 388803:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 388806:4]
  assign ram_opcode_io_deq_bits_MPORT_addr = value_1;
  assign ram_opcode_io_deq_bits_MPORT_data = ram_opcode[ram_opcode_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_opcode_MPORT_data = io_enq_bits_opcode;
  assign ram_opcode_MPORT_addr = value;
  assign ram_opcode_MPORT_mask = 1'h1;
  assign ram_opcode_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_param_io_deq_bits_MPORT_addr = value_1;
  assign ram_param_io_deq_bits_MPORT_data = ram_param[ram_param_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_param_MPORT_data = io_enq_bits_param;
  assign ram_param_MPORT_addr = value;
  assign ram_param_MPORT_mask = 1'h1;
  assign ram_param_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_size_io_deq_bits_MPORT_addr = value_1;
  assign ram_size_io_deq_bits_MPORT_data = ram_size[ram_size_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_size_MPORT_data = io_enq_bits_size;
  assign ram_size_MPORT_addr = value;
  assign ram_size_MPORT_mask = 1'h1;
  assign ram_size_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_source_io_deq_bits_MPORT_addr = value_1;
  assign ram_source_io_deq_bits_MPORT_data = ram_source[ram_source_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_source_MPORT_data = io_enq_bits_source;
  assign ram_source_MPORT_addr = value;
  assign ram_source_MPORT_mask = 1'h1;
  assign ram_source_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_address_io_deq_bits_MPORT_addr = value_1;
  assign ram_address_io_deq_bits_MPORT_data = ram_address[ram_address_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_address_MPORT_data = io_enq_bits_address;
  assign ram_address_MPORT_addr = value;
  assign ram_address_MPORT_mask = 1'h1;
  assign ram_address_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mask_io_deq_bits_MPORT_addr = value_1;
  assign ram_mask_io_deq_bits_MPORT_data = ram_mask[ram_mask_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_mask_MPORT_data = io_enq_bits_mask;
  assign ram_mask_MPORT_addr = value;
  assign ram_mask_MPORT_mask = 1'h1;
  assign ram_mask_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_corrupt_io_deq_bits_MPORT_addr = value_1;
  assign ram_corrupt_io_deq_bits_MPORT_data = ram_corrupt[ram_corrupt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
  assign ram_corrupt_MPORT_data = io_enq_bits_corrupt;
  assign ram_corrupt_MPORT_addr = value;
  assign ram_corrupt_MPORT_mask = 1'h1;
  assign ram_corrupt_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 388812:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 388810:4]
  assign io_deq_bits_opcode = ram_opcode_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388822:4]
  assign io_deq_bits_param = ram_param_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388821:4]
  assign io_deq_bits_size = ram_size_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388820:4]
  assign io_deq_bits_source = ram_source_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388819:4]
  assign io_deq_bits_address = ram_address_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388818:4]
  assign io_deq_bits_mask = ram_mask_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388817:4]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388816:4]
  assign io_deq_bits_corrupt = ram_corrupt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 388815:4]
  always @(posedge clock) begin
    if(ram_opcode_MPORT_en & ram_opcode_MPORT_mask) begin
      ram_opcode[ram_opcode_MPORT_addr] <= ram_opcode_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if(ram_param_MPORT_en & ram_param_MPORT_mask) begin
      ram_param[ram_param_MPORT_addr] <= ram_param_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if(ram_size_MPORT_en & ram_size_MPORT_mask) begin
      ram_size[ram_size_MPORT_addr] <= ram_size_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if(ram_source_MPORT_en & ram_source_MPORT_mask) begin
      ram_source[ram_source_MPORT_addr] <= ram_source_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if(ram_address_MPORT_en & ram_address_MPORT_mask) begin
      ram_address[ram_address_MPORT_addr] <= ram_address_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if(ram_mask_MPORT_en & ram_mask_MPORT_mask) begin
      ram_mask[ram_mask_MPORT_addr] <= ram_mask_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if(ram_corrupt_MPORT_en & ram_corrupt_MPORT_mask) begin
      ram_corrupt[ram_corrupt_MPORT_addr] <= ram_corrupt_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 388771:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388772:4]
      value <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388772:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 388785:4]
      value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 388798:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388773:4]
      value_1 <= 1'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 388773:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 388800:4]
      value_1 <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 388804:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 388774:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 388774:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 388807:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 388808:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[28:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[7:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_corrupt[initvar] = _RAND_7[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  maybe_full = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_20_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 388894:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 388895:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 388896:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [1:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [7:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [1:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [7:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
  input  [63:0] auto_out_d_bits_data // @[chipyard.TestHarness.SmallBoomConfig.fir 388897:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [1:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [7:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [1:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire [7:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [1:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [28:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleOut_0_a_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [1:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [28:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [7:0] bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [7:0] bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
  TLMonitor_55_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 388904:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_44_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388931:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleOut_0_a_q_io_enq_bits_param),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_source(bundleOut_0_a_q_io_enq_bits_source),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleOut_0_a_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_5_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 388945:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 388943:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 388944:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 388957:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 388905:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 388906:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 388943:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 388958:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 388932:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 388933:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388929:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 388946:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 388947:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388929:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388929:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388929:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388929:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 388927:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 388929:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 388902:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 388930:4]
endmodule
module TLMonitor_56_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 388994:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 388995:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 388996:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [2:0]  io_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [2:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [3:0]  io_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [28:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input         io_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [2:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input  [3:0]  io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input         io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 388997:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390488:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390795:4]
  wire  _source_ok_T_4 = io_in_a_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 389014:6]
  wire [12:0] _is_aligned_mask_T_1 = 13'h3f << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 389020:6]
  wire [5:0] is_aligned_mask = ~_is_aligned_mask_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 389022:6]
  wire [28:0] _GEN_71 = {{23'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 389023:6]
  wire [28:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 389023:6]
  wire  is_aligned = _is_aligned_T == 29'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 389024:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 389026:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 389027:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 389029:6]
  wire  _mask_T = io_in_a_bits_size >= 3'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 389030:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 389031:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 389032:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 389033:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389035:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389036:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389038:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389039:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 389040:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 389041:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 389042:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389043:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389044:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389045:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389046:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389047:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389048:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389049:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389050:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389051:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389052:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389053:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389054:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 389055:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 389056:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 389057:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389058:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389059:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389060:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389061:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389062:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389063:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389064:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389065:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389066:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389067:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389068:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389069:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389070:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389071:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389072:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389073:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389074:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389075:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389076:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389077:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389078:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 389079:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 389080:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 389081:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 389088:6]
  wire  _T_20 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 389111:6]
  wire [28:0] _T_33 = io_in_a_bits_address ^ 29'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 389127:8]
  wire [29:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 389128:8]
  wire [29:0] _T_36 = $signed(_T_34) & -30'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 389130:8]
  wire  _T_37 = $signed(_T_36) == 30'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 389131:8]
  wire  _T_43 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389137:8]
  wire  _T_60 = _source_ok_T_4 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389162:8]
  wire  _T_61 = ~_T_60; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389163:8]
  wire  _T_64 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389170:8]
  wire  _T_65 = ~_T_64; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389171:8]
  wire  _T_67 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389177:8]
  wire  _T_68 = ~_T_67; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389178:8]
  wire  _T_69 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 108:27 chipyard.TestHarness.SmallBoomConfig.fir 389183:8]
  wire  _T_71 = _T_69 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389185:8]
  wire  _T_72 = ~_T_71; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389186:8]
  wire [7:0] _T_73 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 389191:8]
  wire  _T_74 = _T_73 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 389192:8]
  wire  _T_76 = _T_74 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389194:8]
  wire  _T_77 = ~_T_76; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389195:8]
  wire  _T_78 = ~io_in_a_bits_corrupt; // @[Monitor.scala 89:18 chipyard.TestHarness.SmallBoomConfig.fir 389200:8]
  wire  _T_80 = _T_78 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389202:8]
  wire  _T_81 = ~_T_80; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389203:8]
  wire  _T_82 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 389209:6]
  wire  _T_135 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 99:31 chipyard.TestHarness.SmallBoomConfig.fir 389289:8]
  wire  _T_137 = _T_135 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389291:8]
  wire  _T_138 = ~_T_137; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389292:8]
  wire  _T_148 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 389315:6]
  wire  _T_164 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 389338:8]
  wire  _T_172 = _T_164 & _T_37; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 389346:8]
  wire  _T_175 = _T_172 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389349:8]
  wire  _T_176 = ~_T_175; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389350:8]
  wire  _T_183 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 109:31 chipyard.TestHarness.SmallBoomConfig.fir 389369:8]
  wire  _T_185 = _T_183 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389371:8]
  wire  _T_186 = ~_T_185; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389372:8]
  wire  _T_187 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 389377:8]
  wire  _T_189 = _T_187 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389379:8]
  wire  _T_190 = ~_T_189; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389380:8]
  wire  _T_195 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 389394:6]
  wire  _T_218 = _source_ok_T_4 & _T_172; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 389420:8]
  wire  _T_220 = _T_218 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389422:8]
  wire  _T_221 = ~_T_220; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389423:8]
  wire  _T_236 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 389459:6]
  wire [7:0] _T_273 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 389515:8]
  wire [7:0] _T_274 = io_in_a_bits_mask & _T_273; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 389516:8]
  wire  _T_275 = _T_274 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 389517:8]
  wire  _T_277 = _T_275 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389519:8]
  wire  _T_278 = ~_T_277; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389520:8]
  wire  _T_279 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 389526:6]
  wire  _T_309 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 138:33 chipyard.TestHarness.SmallBoomConfig.fir 389571:8]
  wire  _T_311 = _T_309 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389573:8]
  wire  _T_312 = ~_T_311; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389574:8]
  wire  _T_317 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 389588:6]
  wire  _T_347 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 145:30 chipyard.TestHarness.SmallBoomConfig.fir 389633:8]
  wire  _T_349 = _T_347 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389635:8]
  wire  _T_350 = ~_T_349; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389636:8]
  wire  _T_355 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 389650:6]
  wire  _T_385 = io_in_a_bits_param <= 3'h1; // @[Bundles.scala 158:28 chipyard.TestHarness.SmallBoomConfig.fir 389695:8]
  wire  _T_387 = _T_385 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389697:8]
  wire  _T_388 = ~_T_387; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389698:8]
  wire  _T_397 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 389722:6]
  wire  _T_399 = _T_397 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389724:6]
  wire  _T_400 = ~_T_399; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389725:6]
  wire  _source_ok_T_10 = io_in_d_bits_source <= 4'h9; // @[Parameters.scala 57:20 chipyard.TestHarness.SmallBoomConfig.fir 389736:6]
  wire  _T_401 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 389742:6]
  wire  _T_403 = _source_ok_T_10 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389745:8]
  wire  _T_404 = ~_T_403; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389746:8]
  wire  _T_405 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 389751:8]
  wire  _T_407 = _T_405 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389753:8]
  wire  _T_408 = ~_T_407; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389754:8]
  wire  _T_409 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 389759:8]
  wire  _T_411 = _T_409 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389761:8]
  wire  _T_412 = ~_T_411; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389762:8]
  wire  _T_413 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 389767:8]
  wire  _T_415 = _T_413 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389769:8]
  wire  _T_416 = ~_T_415; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389770:8]
  wire  _T_417 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 389775:8]
  wire  _T_419 = _T_417 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389777:8]
  wire  _T_420 = ~_T_419; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389778:8]
  wire  _T_421 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 389784:6]
  wire  _T_432 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 389808:8]
  wire  _T_434 = _T_432 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389810:8]
  wire  _T_435 = ~_T_434; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389811:8]
  wire  _T_436 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 389816:8]
  wire  _T_438 = _T_436 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389818:8]
  wire  _T_439 = ~_T_438; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389819:8]
  wire  _T_449 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 389842:6]
  wire  _T_469 = _T_417 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 389883:8]
  wire  _T_471 = _T_469 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389885:8]
  wire  _T_472 = ~_T_471; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389886:8]
  wire  _T_478 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 389901:6]
  wire  _T_495 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 389936:6]
  wire  _T_513 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 389972:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390038:4]
  wire [2:0] a_first_beats1_decode = is_aligned_mask[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 390043:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 390045:4]
  reg [2:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390047:4]
  wire [2:0] a_first_counter1 = a_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390049:4]
  wire  a_first = a_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390050:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 390061:4]
  reg [2:0] param; // @[Monitor.scala 385:22 chipyard.TestHarness.SmallBoomConfig.fir 390062:4]
  reg [2:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 390063:4]
  reg [3:0] source; // @[Monitor.scala 387:22 chipyard.TestHarness.SmallBoomConfig.fir 390064:4]
  reg [28:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 390065:4]
  wire  _T_542 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 390066:4]
  wire  _T_543 = io_in_a_valid & _T_542; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 390067:4]
  wire  _T_544 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 390069:6]
  wire  _T_546 = _T_544 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390071:6]
  wire  _T_547 = ~_T_546; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390072:6]
  wire  _T_548 = io_in_a_bits_param == param; // @[Monitor.scala 391:32 chipyard.TestHarness.SmallBoomConfig.fir 390077:6]
  wire  _T_550 = _T_548 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390079:6]
  wire  _T_551 = ~_T_550; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390080:6]
  wire  _T_552 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 390085:6]
  wire  _T_554 = _T_552 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390087:6]
  wire  _T_555 = ~_T_554; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390088:6]
  wire  _T_556 = io_in_a_bits_source == source; // @[Monitor.scala 393:32 chipyard.TestHarness.SmallBoomConfig.fir 390093:6]
  wire  _T_558 = _T_556 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390095:6]
  wire  _T_559 = ~_T_558; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390096:6]
  wire  _T_560 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 390101:6]
  wire  _T_562 = _T_560 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390103:6]
  wire  _T_563 = ~_T_562; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390104:6]
  wire  _T_565 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 390111:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390119:4]
  wire [12:0] _d_first_beats1_decode_T_1 = 13'h3f << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 390121:4]
  wire [5:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 390123:4]
  wire [2:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[5:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 390124:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 390125:4]
  reg [2:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390127:4]
  wire [2:0] d_first_counter1 = d_first_counter - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390129:4]
  wire  d_first = d_first_counter == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390130:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 390141:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 390142:4]
  reg [2:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 390143:4]
  reg [3:0] source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 390144:4]
  reg  sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 390145:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 390146:4]
  wire  _T_566 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 390147:4]
  wire  _T_567 = io_in_d_valid & _T_566; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 390148:4]
  wire  _T_568 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 390150:6]
  wire  _T_570 = _T_568 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390152:6]
  wire  _T_571 = ~_T_570; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390153:6]
  wire  _T_572 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 390158:6]
  wire  _T_574 = _T_572 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390160:6]
  wire  _T_575 = ~_T_574; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390161:6]
  wire  _T_576 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 390166:6]
  wire  _T_578 = _T_576 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390168:6]
  wire  _T_579 = ~_T_578; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390169:6]
  wire  _T_580 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 390174:6]
  wire  _T_582 = _T_580 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390176:6]
  wire  _T_583 = ~_T_582; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390177:6]
  wire  _T_584 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 390182:6]
  wire  _T_586 = _T_584 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390184:6]
  wire  _T_587 = ~_T_586; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390185:6]
  wire  _T_588 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 390190:6]
  wire  _T_590 = _T_588 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390192:6]
  wire  _T_591 = ~_T_590; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390193:6]
  wire  _T_593 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 390200:4]
  reg [9:0] inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 390209:4]
  reg [39:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 390210:4]
  reg [39:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 390211:4]
  reg [2:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390221:4]
  wire [2:0] a_first_counter1_1 = a_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390223:4]
  wire  a_first_1 = a_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390224:4]
  reg [2:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390243:4]
  wire [2:0] d_first_counter1_1 = d_first_counter_1 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390245:4]
  wire  d_first_1 = d_first_counter_1 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390246:4]
  wire [5:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 390267:4]
  wire [6:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 390267:4]
  wire [39:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 390268:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 390272:4]
  wire [39:0] _GEN_73 = {{24'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 390273:4]
  wire [39:0] _a_opcode_lookup_T_6 = _a_opcode_lookup_T_1 & _GEN_73; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 390273:4]
  wire [39:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[39:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 390274:4]
  wire [39:0] _a_size_lookup_T_1 = inflight_sizes >> _a_opcode_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 390279:4]
  wire [39:0] _a_size_lookup_T_6 = _a_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 390284:4]
  wire [39:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[39:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 390285:4]
  wire  _T_594 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 390309:4]
  wire [15:0] _a_set_wo_ready_T = 16'h1 << io_in_a_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 390312:6]
  wire [15:0] _GEN_15 = _T_594 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 390311:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 390313:6 chipyard.TestHarness.SmallBoomConfig.fir 390260:4]
  wire  _T_597 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 390316:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 390321:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 390322:6]
  wire [3:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 390324:6]
  wire [3:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 4'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 390325:6]
  wire [5:0] _GEN_78 = {io_in_a_bits_source, 2'h0}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 390327:6]
  wire [6:0] _a_opcodes_set_T = {{1'd0}, _GEN_78}; // @[Monitor.scala 656:79 chipyard.TestHarness.SmallBoomConfig.fir 390327:6]
  wire [3:0] a_opcodes_set_interm = _T_597 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390318:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 390323:6 chipyard.TestHarness.SmallBoomConfig.fir 390306:4]
  wire [130:0] _GEN_79 = {{127'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 390328:6]
  wire [130:0] _a_opcodes_set_T_1 = _GEN_79 << _a_opcodes_set_T; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 390328:6]
  wire [3:0] a_sizes_set_interm = _T_597 ? _a_sizes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390318:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 390326:6 chipyard.TestHarness.SmallBoomConfig.fir 390308:4]
  wire [130:0] _GEN_81 = {{127'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 390331:6]
  wire [130:0] _a_sizes_set_T_1 = _GEN_81 << _a_opcodes_set_T; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 390331:6]
  wire [9:0] _T_599 = inflight >> io_in_a_bits_source; // @[Monitor.scala 658:26 chipyard.TestHarness.SmallBoomConfig.fir 390333:6]
  wire  _T_601 = ~_T_599[0]; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 390335:6]
  wire  _T_603 = _T_601 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390337:6]
  wire  _T_604 = ~_T_603; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390338:6]
  wire [15:0] _GEN_16 = _T_597 ? _a_set_wo_ready_T : 16'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390318:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 390320:6 chipyard.TestHarness.SmallBoomConfig.fir 390258:4]
  wire [130:0] _GEN_19 = _T_597 ? _a_opcodes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390318:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 390329:6 chipyard.TestHarness.SmallBoomConfig.fir 390262:4]
  wire [130:0] _GEN_20 = _T_597 ? _a_sizes_set_T_1 : 131'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 390318:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 390332:6 chipyard.TestHarness.SmallBoomConfig.fir 390264:4]
  wire  _T_605 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 390353:4]
  wire  _T_607 = ~_T_401; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 390355:4]
  wire  _T_608 = _T_605 & _T_607; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 390356:4]
  wire [15:0] _d_clr_wo_ready_T = 16'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 390358:6]
  wire [15:0] _GEN_21 = _T_608 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 390357:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 390359:6 chipyard.TestHarness.SmallBoomConfig.fir 390347:4]
  wire  _T_610 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 390362:4]
  wire  _T_613 = _T_610 & _T_607; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 390365:4]
  wire [142:0] _GEN_83 = {{127'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 390374:6]
  wire [142:0] _d_opcodes_clr_T_5 = _GEN_83 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 390374:6]
  wire [15:0] _GEN_22 = _T_613 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 390366:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 390368:6 chipyard.TestHarness.SmallBoomConfig.fir 390345:4]
  wire [142:0] _GEN_23 = _T_613 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 390366:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 390375:6 chipyard.TestHarness.SmallBoomConfig.fir 390349:4]
  wire  _same_cycle_resp_T_2 = io_in_a_bits_source == io_in_d_bits_source; // @[Monitor.scala 681:113 chipyard.TestHarness.SmallBoomConfig.fir 390391:6]
  wire  same_cycle_resp = _T_594 & _same_cycle_resp_T_2; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 390392:6]
  wire [9:0] _T_618 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 390393:6]
  wire  _T_620 = _T_618[0] | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 390395:6]
  wire  _T_622 = _T_620 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390397:6]
  wire  _T_623 = ~_T_622; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390398:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8]
  wire  _T_624 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 390404:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390405:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390405:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390405:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390405:8]
  wire  _T_625 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 390405:8]
  wire  _T_626 = _T_624 | _T_625; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 390406:8]
  wire  _T_628 = _T_626 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390408:8]
  wire  _T_629 = ~_T_628; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390409:8]
  wire  _T_630 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 390414:8]
  wire  _T_632 = _T_630 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390416:8]
  wire  _T_633 = ~_T_632; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390417:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390265:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 390275:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8]
  wire  _T_635 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 390425:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390427:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390427:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390427:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390427:8]
  wire  _T_637 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 390427:8]
  wire  _T_638 = _T_635 | _T_637; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 390428:8]
  wire  _T_640 = _T_638 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390430:8]
  wire  _T_641 = ~_T_640; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390431:8]
  wire [3:0] a_size_lookup = _a_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390276:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 390286:4]
  wire [3:0] _GEN_86 = {{1'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 390436:8]
  wire  _T_642 = _GEN_86 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 390436:8]
  wire  _T_644 = _T_642 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390438:8]
  wire  _T_645 = ~_T_644; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390439:8]
  wire  _T_647 = _T_605 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 390447:4]
  wire  _T_648 = _T_647 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 390448:4]
  wire  _T_650 = _T_648 & _same_cycle_resp_T_2; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 390450:4]
  wire  _T_652 = _T_650 & _T_607; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 390452:4]
  wire  _T_653 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 390454:6]
  wire  _T_654 = _T_653 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 390455:6]
  wire  _T_656 = _T_654 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390457:6]
  wire  _T_657 = ~_T_656; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390458:6]
  wire [9:0] a_set_wo_ready = _GEN_15[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390259:4]
  wire [9:0] d_clr_wo_ready = _GEN_21[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390346:4]
  wire  _T_658 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 390464:4]
  wire  _T_659 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 390465:4]
  wire  _T_660 = ~_T_659; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 390466:4]
  wire  _T_661 = _T_658 | _T_660; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 390467:4]
  wire  _T_663 = _T_661 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390469:4]
  wire  _T_664 = ~_T_663; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390470:4]
  wire [9:0] a_set = _GEN_16[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390257:4]
  wire [9:0] _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 390475:4]
  wire [9:0] d_clr = _GEN_22[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390344:4]
  wire [9:0] _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 390476:4]
  wire [9:0] _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 390477:4]
  wire [39:0] a_opcodes_set = _GEN_19[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390261:4]
  wire [39:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 390479:4]
  wire [39:0] d_opcodes_clr = _GEN_23[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390348:4]
  wire [39:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 390480:4]
  wire [39:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 390481:4]
  wire [39:0] a_sizes_set = _GEN_20[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390263:4]
  wire [39:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 390483:4]
  wire [39:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_opcodes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 390485:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 390487:4]
  wire  _T_665 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 390490:4]
  wire  _T_666 = ~_T_665; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 390491:4]
  wire  _T_667 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 390492:4]
  wire  _T_668 = _T_666 | _T_667; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 390493:4]
  wire  _T_669 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 390494:4]
  wire  _T_670 = _T_668 | _T_669; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 390495:4]
  wire  _T_672 = _T_670 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390497:4]
  wire  _T_673 = ~_T_672; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390498:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 390504:4]
  wire  _T_676 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 390508:4]
  reg [9:0] inflight_1; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 390512:4]
  reg [39:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 390514:4]
  reg [2:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390549:4]
  wire [2:0] d_first_counter1_2 = d_first_counter_2 - 3'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 390551:4]
  wire  d_first_2 = d_first_counter_2 == 3'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 390552:4]
  wire [39:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_opcode_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 390585:4]
  wire [39:0] _c_size_lookup_T_6 = _c_size_lookup_T_1 & _GEN_73; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 390590:4]
  wire [39:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[39:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 390591:4]
  wire  _T_694 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 390669:4]
  wire  _T_696 = _T_694 & _T_401; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 390671:4]
  wire  _T_698 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 390677:4]
  wire  _T_700 = _T_698 & _T_401; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 390679:4]
  wire [15:0] _GEN_67 = _T_700 ? _d_clr_wo_ready_T : 16'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 390680:4 Monitor.scala 784:21 chipyard.TestHarness.SmallBoomConfig.fir 390682:6 chipyard.TestHarness.SmallBoomConfig.fir 390661:4]
  wire [142:0] _GEN_68 = _T_700 ? _d_opcodes_clr_T_5 : 143'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 390680:4 Monitor.scala 785:21 chipyard.TestHarness.SmallBoomConfig.fir 390689:6 chipyard.TestHarness.SmallBoomConfig.fir 390665:4]
  wire [9:0] _T_704 = inflight_1 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 390715:6]
  wire  _T_708 = _T_704[0] | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390719:6]
  wire  _T_709 = ~_T_708; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390720:6]
  wire [3:0] c_size_lookup = _c_size_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390573:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 390592:4]
  wire  _T_714 = _GEN_86 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 390738:8]
  wire  _T_716 = _T_714 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390740:8]
  wire  _T_717 = ~_T_716; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390741:8]
  wire [9:0] d_clr_1 = _GEN_67[9:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390660:4]
  wire [9:0] _inflight_T_4 = ~d_clr_1; // @[Monitor.scala 809:46 chipyard.TestHarness.SmallBoomConfig.fir 390783:4]
  wire [9:0] _inflight_T_5 = inflight_1 & _inflight_T_4; // @[Monitor.scala 809:44 chipyard.TestHarness.SmallBoomConfig.fir 390784:4]
  wire [39:0] d_opcodes_clr_1 = _GEN_68[39:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 390664:4]
  wire [39:0] _inflight_opcodes_T_4 = ~d_opcodes_clr_1; // @[Monitor.scala 810:62 chipyard.TestHarness.SmallBoomConfig.fir 390787:4]
  wire [39:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_opcodes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 390792:4]
  reg [31:0] watchdog_1; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 390794:4]
  wire  _T_734 = |inflight_1; // @[Monitor.scala 816:26 chipyard.TestHarness.SmallBoomConfig.fir 390797:4]
  wire  _T_735 = ~_T_734; // @[Monitor.scala 816:16 chipyard.TestHarness.SmallBoomConfig.fir 390798:4]
  wire  _T_736 = plusarg_reader_1_out == 32'h0; // @[Monitor.scala 816:39 chipyard.TestHarness.SmallBoomConfig.fir 390799:4]
  wire  _T_737 = _T_735 | _T_736; // @[Monitor.scala 816:30 chipyard.TestHarness.SmallBoomConfig.fir 390800:4]
  wire  _T_738 = watchdog_1 < plusarg_reader_1_out; // @[Monitor.scala 816:59 chipyard.TestHarness.SmallBoomConfig.fir 390801:4]
  wire  _T_739 = _T_737 | _T_738; // @[Monitor.scala 816:47 chipyard.TestHarness.SmallBoomConfig.fir 390802:4]
  wire  _T_741 = _T_739 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390804:4]
  wire  _T_742 = ~_T_741; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390805:4]
  wire [31:0] _watchdog_T_3 = watchdog_1 + 32'h1; // @[Monitor.scala 818:26 chipyard.TestHarness.SmallBoomConfig.fir 390811:4]
  wire  _GEN_98 = io_in_a_valid & _T_20; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389139:10]
  wire  _GEN_114 = io_in_a_valid & _T_82; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389237:10]
  wire  _GEN_132 = io_in_a_valid & _T_148; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389334:10]
  wire  _GEN_146 = io_in_a_valid & _T_195; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389425:10]
  wire  _GEN_156 = io_in_a_valid & _T_236; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389490:10]
  wire  _GEN_166 = io_in_a_valid & _T_279; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389554:10]
  wire  _GEN_176 = io_in_a_valid & _T_317; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389616:10]
  wire  _GEN_186 = io_in_a_valid & _T_355; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389678:10]
  wire  _GEN_198 = io_in_d_valid & _T_401; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389748:10]
  wire  _GEN_208 = io_in_d_valid & _T_421; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389790:10]
  wire  _GEN_222 = io_in_d_valid & _T_449; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389848:10]
  wire  _GEN_236 = io_in_d_valid & _T_478; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389907:10]
  wire  _GEN_244 = io_in_d_valid & _T_495; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389942:10]
  wire  _GEN_252 = io_in_d_valid & _T_513; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389978:10]
  wire  _GEN_260 = _T_608 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390411:10]
  wire  _GEN_265 = _T_608 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390433:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390488:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 390795:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390047:4]
      a_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390047:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390057:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390058:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390046:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 3'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390112:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 390113:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390112:4]
      param <= io_in_a_bits_param; // @[Monitor.scala 398:15 chipyard.TestHarness.SmallBoomConfig.fir 390114:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390112:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 390115:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390112:4]
      source <= io_in_a_bits_source; // @[Monitor.scala 400:15 chipyard.TestHarness.SmallBoomConfig.fir 390116:6]
    end
    if (_T_565) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 390112:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 390117:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390127:4]
      d_first_counter <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390127:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390137:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390138:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390126:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 3'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390201:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 390202:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390201:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 390203:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390201:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 390204:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390201:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 390205:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390201:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 390206:6]
    end
    if (_T_593) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 390201:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 390207:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 390209:4]
      inflight <= 10'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 390209:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 390478:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 390210:4]
      inflight_opcodes <= 40'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 390210:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 390482:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 390211:4]
      inflight_sizes <= 40'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 390211:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 390486:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390221:4]
      a_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390221:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390231:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390232:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390046:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 3'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390243:4]
      d_first_counter_1 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390243:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390253:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390254:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390126:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 3'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 390487:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 390487:4]
    end else if (_T_676) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 390509:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 390510:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 390505:4]
    end
    if (reset) begin // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 390512:4]
      inflight_1 <= 10'h0; // @[Monitor.scala 723:35 chipyard.TestHarness.SmallBoomConfig.fir 390512:4]
    end else begin
      inflight_1 <= _inflight_T_5; // @[Monitor.scala 809:22 chipyard.TestHarness.SmallBoomConfig.fir 390785:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 390514:4]
      inflight_sizes_1 <= 40'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 390514:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 390793:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390549:4]
      d_first_counter_2 <= 3'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 390549:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 390559:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 390560:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 390126:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 3'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    if (reset) begin // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 390794:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 813:27 chipyard.TestHarness.SmallBoomConfig.fir 390794:4]
    end else if (_d_first_T) begin // @[Monitor.scala 819:47 chipyard.TestHarness.SmallBoomConfig.fir 390818:4]
      watchdog_1 <= 32'h0; // @[Monitor.scala 819:58 chipyard.TestHarness.SmallBoomConfig.fir 390819:6]
    end else begin
      watchdog_1 <= _watchdog_T_3; // @[Monitor.scala 818:14 chipyard.TestHarness.SmallBoomConfig.fir 390812:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_20 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389139:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389140:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389158:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389159:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389165:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389166:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389173:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389174:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389180:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389181:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389188:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389189:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389197:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389198:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389205:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_98 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389206:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_82 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389237:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389238:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389256:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389257:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389263:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389264:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389271:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_65) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389272:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389278:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389279:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389286:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_72) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389287:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389294:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_138) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389295:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389303:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_77) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389304:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389311:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_114 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389312:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_148 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389334:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389335:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389352:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_176) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389353:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389359:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389360:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389366:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389367:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389374:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389375:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389382:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389383:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389390:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389391:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_195 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389425:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389426:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389432:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389433:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389439:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389440:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389447:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389448:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389455:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_146 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389456:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_236 & _T_221) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389490:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_221) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389491:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389497:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389498:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389504:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389505:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389512:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_186) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389513:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389522:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_156 & _T_278) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389523:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_279 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389554:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389555:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389561:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389562:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389568:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389569:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389576:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_312) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389577:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389584:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_166 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389585:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_317 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389616:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389617:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389623:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389624:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389630:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389631:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389638:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_350) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389639:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389646:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_176 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389647:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_355 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389678:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_43) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389679:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389685:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_61) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389686:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389692:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_68) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389693:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint carries invalid opcode param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389700:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_388) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389701:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389708:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_190) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389709:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389716:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_81) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 389717:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389727:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_400) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389728:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_401 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389748:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389749:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389756:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389757:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389764:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389765:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389772:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389773:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389780:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389781:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_421 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389790:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389791:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389797:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389798:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389805:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389806:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389813:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389814:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389821:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389822:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389829:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389830:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389838:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_208 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389839:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_449 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389848:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389849:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389855:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_43) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389856:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389863:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_408) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389864:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389871:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_435) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389872:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389879:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_439) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389880:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389888:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389889:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389897:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_222 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389898:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_478 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389907:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389908:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389915:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389916:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389923:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389924:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389932:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_236 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389933:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_495 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389942:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389943:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389950:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389951:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389959:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_472) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389960:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389968:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_244 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389969:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_513 & _T_404) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389978:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_404) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389979:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389986:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_412) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389987:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389994:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_416) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 389995:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is denied (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390003:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_252 & _T_420) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390004:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390074:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_547) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390075:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390082:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_551) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390083:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390090:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_555) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390091:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390098:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_559) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390099:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390106:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_543 & _T_563) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390107:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390155:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_571) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390156:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390163:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_575) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390164:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390171:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_579) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390172:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390179:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_583) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390180:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390187:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_587) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390188:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390195:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_567 & _T_591) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390196:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390340:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597 & _T_604) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390341:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390400:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_608 & _T_623) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390401:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & same_cycle_resp & _T_629) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390411:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_629) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390412:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390419:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_260 & _T_633) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390420:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_608 & ~same_cycle_resp & _T_641) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390433:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_641) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390434:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390441:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_265 & _T_645) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390442:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390460:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_652 & _T_657) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390461:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_664) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390472:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_664) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390473:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_673) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390500:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_673) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390501:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390722:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_709) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390723:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390743:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_696 & _T_717) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 390744:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:328:92)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390807:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 390808:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  d_first_counter = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  opcode_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  param_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  size_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  source_1 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  sink = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  denied = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inflight = _RAND_13[9:0];
  _RAND_14 = {2{`RANDOM}};
  inflight_opcodes = _RAND_14[39:0];
  _RAND_15 = {2{`RANDOM}};
  inflight_sizes = _RAND_15[39:0];
  _RAND_16 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  watchdog = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inflight_1 = _RAND_19[9:0];
  _RAND_20 = {2{`RANDOM}};
  inflight_sizes_1 = _RAND_20[39:0];
  _RAND_21 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  watchdog_1 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater_7_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 390822:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 390823:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 390824:4]
  input         io_repeat, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output        io_full, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output        io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input         io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input  [2:0]  io_enq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input  [2:0]  io_enq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input  [2:0]  io_enq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input  [3:0]  io_enq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input  [28:0] io_enq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input  [7:0]  io_enq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input         io_enq_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  input         io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output        io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output [2:0]  io_deq_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output [2:0]  io_deq_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output [2:0]  io_deq_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output [3:0]  io_deq_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output [28:0] io_deq_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output [7:0]  io_deq_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
  output        io_deq_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 390825:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390827:4]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390828:4]
  reg [2:0] saved_param; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390828:4]
  reg [2:0] saved_size; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390828:4]
  reg [3:0] saved_source; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390828:4]
  reg [28:0] saved_address; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390828:4]
  reg [7:0] saved_mask; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390828:4]
  reg  saved_corrupt; // @[Repeater.scala 20:18 chipyard.TestHarness.SmallBoomConfig.fir 390828:4]
  wire  _io_enq_ready_T = ~full; // @[Repeater.scala 24:35 chipyard.TestHarness.SmallBoomConfig.fir 390831:4]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390844:4]
  wire  _T_1 = _T & io_repeat; // @[Repeater.scala 28:23 chipyard.TestHarness.SmallBoomConfig.fir 390845:4]
  wire  _GEN_0 = _T_1 | full; // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4 Repeater.scala 28:45 chipyard.TestHarness.SmallBoomConfig.fir 390847:6 Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390827:4]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390857:4]
  wire  _T_3 = ~io_repeat; // @[Repeater.scala 29:26 chipyard.TestHarness.SmallBoomConfig.fir 390858:4]
  wire  _T_4 = _T_2 & _T_3; // @[Repeater.scala 29:23 chipyard.TestHarness.SmallBoomConfig.fir 390859:4]
  assign io_full = full; // @[Repeater.scala 26:11 chipyard.TestHarness.SmallBoomConfig.fir 390843:4]
  assign io_enq_ready = io_deq_ready & _io_enq_ready_T; // @[Repeater.scala 24:32 chipyard.TestHarness.SmallBoomConfig.fir 390832:4]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32 chipyard.TestHarness.SmallBoomConfig.fir 390829:4]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390834:4]
  assign io_deq_bits_param = full ? saved_param : io_enq_bits_param; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390834:4]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390834:4]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390834:4]
  assign io_deq_bits_address = full ? saved_address : io_enq_bits_address; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390834:4]
  assign io_deq_bits_mask = full ? saved_mask : io_enq_bits_mask; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390834:4]
  assign io_deq_bits_corrupt = full ? saved_corrupt : io_enq_bits_corrupt; // @[Repeater.scala 25:21 chipyard.TestHarness.SmallBoomConfig.fir 390834:4]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390827:4]
      full <= 1'h0; // @[Repeater.scala 19:21 chipyard.TestHarness.SmallBoomConfig.fir 390827:4]
    end else if (_T_4) begin // @[Repeater.scala 29:38 chipyard.TestHarness.SmallBoomConfig.fir 390860:4]
      full <= 1'h0; // @[Repeater.scala 29:45 chipyard.TestHarness.SmallBoomConfig.fir 390861:6]
    end else begin
      full <= _GEN_0;
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390855:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
      saved_param <= io_enq_bits_param; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390854:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390853:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390852:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
      saved_address <= io_enq_bits_address; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390851:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
      saved_mask <= io_enq_bits_mask; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390850:6]
    end
    if (_T_1) begin // @[Repeater.scala 28:38 chipyard.TestHarness.SmallBoomConfig.fir 390846:4]
      saved_corrupt <= io_enq_bits_corrupt; // @[Repeater.scala 28:62 chipyard.TestHarness.SmallBoomConfig.fir 390848:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  saved_source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  saved_address = _RAND_5[28:0];
  _RAND_6 = {1{`RANDOM}};
  saved_mask = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  saved_corrupt = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLFragmenter_7_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 390864:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 390865:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 390866:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [2:0]  auto_in_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [2:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [3:0]  auto_in_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [28:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_in_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [2:0]  auto_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [1:0]  auto_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [2:0]  auto_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [3:0]  auto_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output        auto_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output        auto_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output        auto_in_d_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [1:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [7:0]  auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [28:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [1:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [7:0]  auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 390867:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [2:0] monitor_io_in_a_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [2:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [3:0] monitor_io_in_a_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [28:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_a_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [2:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire [3:0] monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
  wire  repeater_clock; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_reset; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_repeat; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_full; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_enq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_enq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [2:0] repeater_io_enq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [2:0] repeater_io_enq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [2:0] repeater_io_enq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [3:0] repeater_io_enq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [28:0] repeater_io_enq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [7:0] repeater_io_enq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_enq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_deq_ready; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_deq_valid; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [2:0] repeater_io_deq_bits_opcode; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [2:0] repeater_io_deq_bits_param; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [2:0] repeater_io_deq_bits_size; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [3:0] repeater_io_deq_bits_source; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [28:0] repeater_io_deq_bits_address; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire [7:0] repeater_io_deq_bits_mask; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  wire  repeater_io_deq_bits_corrupt; // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
  reg [2:0] acknum; // @[Fragmenter.scala 189:29 chipyard.TestHarness.SmallBoomConfig.fir 390901:4]
  reg [2:0] dOrig; // @[Fragmenter.scala 190:24 chipyard.TestHarness.SmallBoomConfig.fir 390902:4]
  reg  dToggle; // @[Fragmenter.scala 191:30 chipyard.TestHarness.SmallBoomConfig.fir 390903:4]
  wire [2:0] dFragnum = auto_out_d_bits_source[2:0]; // @[Fragmenter.scala 192:41 chipyard.TestHarness.SmallBoomConfig.fir 390904:4]
  wire  dFirst = acknum == 3'h0; // @[Fragmenter.scala 193:29 chipyard.TestHarness.SmallBoomConfig.fir 390905:4]
  wire  dLast = dFragnum == 3'h0; // @[Fragmenter.scala 194:30 chipyard.TestHarness.SmallBoomConfig.fir 390906:4]
  wire [3:0] dsizeOH = 4'h1 << auto_out_d_bits_size; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 390908:4]
  wire [5:0] _dsizeOH1_T_1 = 6'h7 << auto_out_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 390911:4]
  wire [2:0] dsizeOH1 = ~_dsizeOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 390913:4]
  wire  dHasData = auto_out_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 390914:4]
  wire  ack_decrement = dHasData | dsizeOH[3]; // @[Fragmenter.scala 204:32 chipyard.TestHarness.SmallBoomConfig.fir 390931:4]
  wire [5:0] _dFirst_size_T = {dFragnum, 3'h0}; // @[Fragmenter.scala 206:47 chipyard.TestHarness.SmallBoomConfig.fir 390932:4]
  wire [5:0] _GEN_7 = {{3'd0}, dsizeOH1}; // @[Fragmenter.scala 206:69 chipyard.TestHarness.SmallBoomConfig.fir 390933:4]
  wire [5:0] dFirst_size_lo = _dFirst_size_T | _GEN_7; // @[Fragmenter.scala 206:69 chipyard.TestHarness.SmallBoomConfig.fir 390933:4]
  wire [6:0] _dFirst_size_T_1 = {dFirst_size_lo, 1'h0}; // @[package.scala 232:35 chipyard.TestHarness.SmallBoomConfig.fir 390934:4]
  wire [6:0] _dFirst_size_T_2 = _dFirst_size_T_1 | 7'h1; // @[package.scala 232:40 chipyard.TestHarness.SmallBoomConfig.fir 390935:4]
  wire [6:0] _dFirst_size_T_3 = {1'h0,dFirst_size_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 390936:4]
  wire [6:0] _dFirst_size_T_4 = ~_dFirst_size_T_3; // @[package.scala 232:53 chipyard.TestHarness.SmallBoomConfig.fir 390937:4]
  wire [6:0] _dFirst_size_T_5 = _dFirst_size_T_2 & _dFirst_size_T_4; // @[package.scala 232:51 chipyard.TestHarness.SmallBoomConfig.fir 390938:4]
  wire [2:0] dFirst_size_hi = _dFirst_size_T_5[6:4]; // @[OneHot.scala 30:18 chipyard.TestHarness.SmallBoomConfig.fir 390939:4]
  wire [3:0] dFirst_size_lo_1 = _dFirst_size_T_5[3:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.SmallBoomConfig.fir 390940:4]
  wire  dFirst_size_hi_1 = |dFirst_size_hi; // @[OneHot.scala 32:14 chipyard.TestHarness.SmallBoomConfig.fir 390941:4]
  wire [3:0] _GEN_8 = {{1'd0}, dFirst_size_hi}; // @[OneHot.scala 32:28 chipyard.TestHarness.SmallBoomConfig.fir 390942:4]
  wire [3:0] _dFirst_size_T_6 = _GEN_8 | dFirst_size_lo_1; // @[OneHot.scala 32:28 chipyard.TestHarness.SmallBoomConfig.fir 390942:4]
  wire [1:0] dFirst_size_hi_2 = _dFirst_size_T_6[3:2]; // @[OneHot.scala 30:18 chipyard.TestHarness.SmallBoomConfig.fir 390943:4]
  wire [1:0] dFirst_size_lo_2 = _dFirst_size_T_6[1:0]; // @[OneHot.scala 31:18 chipyard.TestHarness.SmallBoomConfig.fir 390944:4]
  wire  dFirst_size_hi_3 = |dFirst_size_hi_2; // @[OneHot.scala 32:14 chipyard.TestHarness.SmallBoomConfig.fir 390945:4]
  wire [1:0] _dFirst_size_T_7 = dFirst_size_hi_2 | dFirst_size_lo_2; // @[OneHot.scala 32:28 chipyard.TestHarness.SmallBoomConfig.fir 390946:4]
  wire  dFirst_size_lo_3 = _dFirst_size_T_7[1]; // @[CircuitMath.scala 30:8 chipyard.TestHarness.SmallBoomConfig.fir 390947:4]
  wire [2:0] dFirst_size = {dFirst_size_hi_1,dFirst_size_hi_3,dFirst_size_lo_3}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 390949:4]
  wire  _drop_T = ~dHasData; // @[Fragmenter.scala 222:20 chipyard.TestHarness.SmallBoomConfig.fir 390962:4]
  wire  _drop_T_2 = ~dLast; // @[Fragmenter.scala 222:33 chipyard.TestHarness.SmallBoomConfig.fir 390964:4]
  wire  drop = _drop_T & _drop_T_2; // @[Fragmenter.scala 222:30 chipyard.TestHarness.SmallBoomConfig.fir 390965:4]
  wire  bundleOut_0_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.SmallBoomConfig.fir 390966:4]
  wire  _T_7 = bundleOut_0_d_ready & auto_out_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 390950:4]
  wire [2:0] _GEN_9 = {{2'd0}, ack_decrement}; // @[Fragmenter.scala 209:55 chipyard.TestHarness.SmallBoomConfig.fir 390952:6]
  wire [2:0] _acknum_T_1 = acknum - _GEN_9; // @[Fragmenter.scala 209:55 chipyard.TestHarness.SmallBoomConfig.fir 390953:6]
  wire  _bundleIn_0_d_valid_T = ~drop; // @[Fragmenter.scala 224:39 chipyard.TestHarness.SmallBoomConfig.fir 390968:4]
  wire  _aFrag_T = repeater_io_deq_bits_size > 3'h3; // @[Fragmenter.scala 285:31 chipyard.TestHarness.SmallBoomConfig.fir 391001:4]
  wire [2:0] aFrag = _aFrag_T ? 3'h3 : repeater_io_deq_bits_size; // @[Fragmenter.scala 285:24 chipyard.TestHarness.SmallBoomConfig.fir 391002:4]
  wire [12:0] _aOrigOH1_T_1 = 13'h3f << repeater_io_deq_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 391004:4]
  wire [5:0] aOrigOH1 = ~_aOrigOH1_T_1[5:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 391006:4]
  wire [9:0] _aFragOH1_T_1 = 10'h7 << aFrag; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 391008:4]
  wire [2:0] aFragOH1 = ~_aFragOH1_T_1[2:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 391010:4]
  wire  aHasData = ~repeater_io_deq_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 391012:4]
  reg [2:0] gennum; // @[Fragmenter.scala 291:29 chipyard.TestHarness.SmallBoomConfig.fir 391014:4]
  wire  aFirst = gennum == 3'h0; // @[Fragmenter.scala 292:29 chipyard.TestHarness.SmallBoomConfig.fir 391015:4]
  wire [2:0] _old_gennum1_T_2 = gennum - 3'h1; // @[Fragmenter.scala 293:79 chipyard.TestHarness.SmallBoomConfig.fir 391018:4]
  wire [2:0] old_gennum1 = aFirst ? aOrigOH1[5:3] : _old_gennum1_T_2; // @[Fragmenter.scala 293:30 chipyard.TestHarness.SmallBoomConfig.fir 391019:4]
  wire [2:0] _new_gennum_T = ~old_gennum1; // @[Fragmenter.scala 294:28 chipyard.TestHarness.SmallBoomConfig.fir 391020:4]
  wire [2:0] new_gennum = ~_new_gennum_T; // @[Fragmenter.scala 294:26 chipyard.TestHarness.SmallBoomConfig.fir 391023:4]
  reg  aToggle_r; // @[Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 391030:4]
  wire  _GEN_5 = aFirst ? dToggle : aToggle_r; // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 391031:4 Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 391032:6 Reg.scala 15:16 chipyard.TestHarness.SmallBoomConfig.fir 391030:4]
  wire  bundleOut_0_a_bits_source_hi_lo = ~_GEN_5; // @[Fragmenter.scala 297:23 chipyard.TestHarness.SmallBoomConfig.fir 391035:4]
  wire  bundleOut_0_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391044:4]
  wire  _T_8 = auto_out_a_ready & bundleOut_0_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 391036:4]
  wire  _repeater_io_repeat_T = ~aHasData; // @[Fragmenter.scala 302:31 chipyard.TestHarness.SmallBoomConfig.fir 391040:4]
  wire  _repeater_io_repeat_T_1 = new_gennum != 3'h0; // @[Fragmenter.scala 302:53 chipyard.TestHarness.SmallBoomConfig.fir 391041:4]
  wire [5:0] _bundleOut_0_a_bits_address_T = {old_gennum1, 3'h0}; // @[Fragmenter.scala 304:65 chipyard.TestHarness.SmallBoomConfig.fir 391045:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_1 = ~aOrigOH1; // @[Fragmenter.scala 304:90 chipyard.TestHarness.SmallBoomConfig.fir 391046:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_2 = _bundleOut_0_a_bits_address_T | _bundleOut_0_a_bits_address_T_1; // @[Fragmenter.scala 304:88 chipyard.TestHarness.SmallBoomConfig.fir 391047:4]
  wire [5:0] _GEN_10 = {{3'd0}, aFragOH1}; // @[Fragmenter.scala 304:100 chipyard.TestHarness.SmallBoomConfig.fir 391048:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_3 = _bundleOut_0_a_bits_address_T_2 | _GEN_10; // @[Fragmenter.scala 304:100 chipyard.TestHarness.SmallBoomConfig.fir 391048:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_4 = _bundleOut_0_a_bits_address_T_3 | 6'h7; // @[Fragmenter.scala 304:111 chipyard.TestHarness.SmallBoomConfig.fir 391049:4]
  wire [5:0] _bundleOut_0_a_bits_address_T_5 = ~_bundleOut_0_a_bits_address_T_4; // @[Fragmenter.scala 304:51 chipyard.TestHarness.SmallBoomConfig.fir 391050:4]
  wire [28:0] _GEN_11 = {{23'd0}, _bundleOut_0_a_bits_address_T_5}; // @[Fragmenter.scala 304:49 chipyard.TestHarness.SmallBoomConfig.fir 391051:4]
  wire [4:0] bundleOut_0_a_bits_source_hi = {repeater_io_deq_bits_source,bundleOut_0_a_bits_source_hi_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 391053:4]
  wire  _T_9 = ~repeater_io_full; // @[Fragmenter.scala 309:17 chipyard.TestHarness.SmallBoomConfig.fir 391057:4]
  wire  _T_11 = _T_9 | _repeater_io_repeat_T; // @[Fragmenter.scala 309:35 chipyard.TestHarness.SmallBoomConfig.fir 391059:4]
  wire  _T_13 = _T_11 | reset; // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391061:4]
  wire  _T_14 = ~_T_13; // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391062:4]
  wire  _T_16 = repeater_io_deq_bits_mask == 8'hff; // @[Fragmenter.scala 312:53 chipyard.TestHarness.SmallBoomConfig.fir 391069:4]
  wire  _T_17 = _T_9 | _T_16; // @[Fragmenter.scala 312:35 chipyard.TestHarness.SmallBoomConfig.fir 391070:4]
  wire  _T_19 = _T_17 | reset; // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391072:4]
  wire  _T_20 = ~_T_19; // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391073:4]
  TLMonitor_56_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 390874:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(monitor_io_in_a_bits_param),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_source(monitor_io_in_a_bits_source),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(monitor_io_in_a_bits_corrupt),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Repeater_7_inTestHarness repeater ( // @[Fragmenter.scala 262:30 chipyard.TestHarness.SmallBoomConfig.fir 390976:4]
    .clock(repeater_clock),
    .reset(repeater_reset),
    .io_repeat(repeater_io_repeat),
    .io_full(repeater_io_full),
    .io_enq_ready(repeater_io_enq_ready),
    .io_enq_valid(repeater_io_enq_valid),
    .io_enq_bits_opcode(repeater_io_enq_bits_opcode),
    .io_enq_bits_param(repeater_io_enq_bits_param),
    .io_enq_bits_size(repeater_io_enq_bits_size),
    .io_enq_bits_source(repeater_io_enq_bits_source),
    .io_enq_bits_address(repeater_io_enq_bits_address),
    .io_enq_bits_mask(repeater_io_enq_bits_mask),
    .io_enq_bits_corrupt(repeater_io_enq_bits_corrupt),
    .io_deq_ready(repeater_io_deq_ready),
    .io_deq_valid(repeater_io_deq_valid),
    .io_deq_bits_opcode(repeater_io_deq_bits_opcode),
    .io_deq_bits_param(repeater_io_deq_bits_param),
    .io_deq_bits_size(repeater_io_deq_bits_size),
    .io_deq_bits_source(repeater_io_deq_bits_source),
    .io_deq_bits_address(repeater_io_deq_bits_address),
    .io_deq_bits_mask(repeater_io_deq_bits_mask),
    .io_deq_bits_corrupt(repeater_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 Fragmenter.scala 263:25 chipyard.TestHarness.SmallBoomConfig.fir 390980:4]
  assign auto_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.SmallBoomConfig.fir 390969:4]
  assign auto_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign auto_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign auto_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.SmallBoomConfig.fir 390974:4]
  assign auto_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.SmallBoomConfig.fir 390972:4]
  assign auto_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign auto_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign auto_in_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign auto_out_a_valid = repeater_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391044:4]
  assign auto_out_a_bits_opcode = repeater_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391044:4]
  assign auto_out_a_bits_param = repeater_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391044:4]
  assign auto_out_a_bits_size = aFrag[1:0]; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 Fragmenter.scala 306:25 chipyard.TestHarness.SmallBoomConfig.fir 391056:4]
  assign auto_out_a_bits_source = {bundleOut_0_a_bits_source_hi,new_gennum}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 391054:4]
  assign auto_out_a_bits_address = repeater_io_deq_bits_address | _GEN_11; // @[Fragmenter.scala 304:49 chipyard.TestHarness.SmallBoomConfig.fir 391051:4]
  assign auto_out_a_bits_mask = repeater_io_full ? 8'hff : auto_in_a_bits_mask; // @[Fragmenter.scala 313:31 chipyard.TestHarness.SmallBoomConfig.fir 391078:4]
  assign auto_out_a_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign auto_out_a_bits_corrupt = repeater_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 Fragmenter.scala 303:15 chipyard.TestHarness.SmallBoomConfig.fir 391044:4]
  assign auto_out_d_ready = auto_in_d_ready | drop; // @[Fragmenter.scala 223:35 chipyard.TestHarness.SmallBoomConfig.fir 390966:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 390875:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 390876:4]
  assign monitor_io_in_a_ready = repeater_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 Fragmenter.scala 263:25 chipyard.TestHarness.SmallBoomConfig.fir 390980:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign monitor_io_in_d_valid = auto_out_d_valid & _bundleIn_0_d_valid_T; // @[Fragmenter.scala 224:36 chipyard.TestHarness.SmallBoomConfig.fir 390969:4]
  assign monitor_io_in_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign monitor_io_in_d_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign monitor_io_in_d_bits_size = dFirst ? dFirst_size : dOrig; // @[Fragmenter.scala 227:32 chipyard.TestHarness.SmallBoomConfig.fir 390974:4]
  assign monitor_io_in_d_bits_source = auto_out_d_bits_source[7:4]; // @[Fragmenter.scala 226:47 chipyard.TestHarness.SmallBoomConfig.fir 390972:4]
  assign monitor_io_in_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign monitor_io_in_d_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign monitor_io_in_d_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  assign repeater_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 390978:4]
  assign repeater_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 390979:4]
  assign repeater_io_repeat = _repeater_io_repeat_T & _repeater_io_repeat_T_1; // @[Fragmenter.scala 302:41 chipyard.TestHarness.SmallBoomConfig.fir 391042:4]
  assign repeater_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_enq_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_enq_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_enq_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 390872:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 390900:4]
  assign repeater_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 390897:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 390899:4]
  always @(posedge clock) begin
    if (reset) begin // @[Fragmenter.scala 189:29 chipyard.TestHarness.SmallBoomConfig.fir 390901:4]
      acknum <= 3'h0; // @[Fragmenter.scala 189:29 chipyard.TestHarness.SmallBoomConfig.fir 390901:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.SmallBoomConfig.fir 390951:4]
      if (dFirst) begin // @[Fragmenter.scala 209:24 chipyard.TestHarness.SmallBoomConfig.fir 390954:6]
        acknum <= dFragnum;
      end else begin
        acknum <= _acknum_T_1;
      end
    end
    if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.SmallBoomConfig.fir 390951:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.SmallBoomConfig.fir 390956:6]
        dOrig <= dFirst_size; // @[Fragmenter.scala 211:19 chipyard.TestHarness.SmallBoomConfig.fir 390957:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 191:30 chipyard.TestHarness.SmallBoomConfig.fir 390903:4]
      dToggle <= 1'h0; // @[Fragmenter.scala 191:30 chipyard.TestHarness.SmallBoomConfig.fir 390903:4]
    end else if (_T_7) begin // @[Fragmenter.scala 208:29 chipyard.TestHarness.SmallBoomConfig.fir 390951:4]
      if (dFirst) begin // @[Fragmenter.scala 210:25 chipyard.TestHarness.SmallBoomConfig.fir 390956:6]
        dToggle <= auto_out_d_bits_source[3]; // @[Fragmenter.scala 212:21 chipyard.TestHarness.SmallBoomConfig.fir 390959:8]
      end
    end
    if (reset) begin // @[Fragmenter.scala 291:29 chipyard.TestHarness.SmallBoomConfig.fir 391014:4]
      gennum <= 3'h0; // @[Fragmenter.scala 291:29 chipyard.TestHarness.SmallBoomConfig.fir 391014:4]
    end else if (_T_8) begin // @[Fragmenter.scala 300:29 chipyard.TestHarness.SmallBoomConfig.fir 391037:4]
      gennum <= new_gennum; // @[Fragmenter.scala 300:38 chipyard.TestHarness.SmallBoomConfig.fir 391038:6]
    end
    if (aFirst) begin // @[Reg.scala 16:19 chipyard.TestHarness.SmallBoomConfig.fir 391031:4]
      aToggle_r <= dToggle; // @[Reg.scala 16:23 chipyard.TestHarness.SmallBoomConfig.fir 391032:6]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_14) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:309 assert (!repeater.io.full || !aHasData)\n"
            ); // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391064:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_14) begin
          $fatal; // @[Fragmenter.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 391065:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Fragmenter.scala:312 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n"
            ); // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391075:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_20) begin
          $fatal; // @[Fragmenter.scala 312:16 chipyard.TestHarness.SmallBoomConfig.fir 391076:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  acknum = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dOrig = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  gennum = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  aToggle_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLMonitor_57_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 391116:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 391117:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 391118:4]
  input         io_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input         io_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [2:0]  io_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [3:0]  io_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [31:0] io_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [7:0]  io_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input         io_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input         io_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [2:0]  io_in_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [1:0]  io_in_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [3:0]  io_in_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input         io_in_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input  [2:0]  io_in_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input         io_in_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
  input         io_in_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 391119:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393058:4]
  wire [31:0] plusarg_reader_1_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393365:4]
  wire [26:0] _is_aligned_mask_T_1 = 27'hfff << io_in_a_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 391135:6]
  wire [11:0] is_aligned_mask = ~_is_aligned_mask_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 391137:6]
  wire [31:0] _GEN_71 = {{20'd0}, is_aligned_mask}; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 391138:6]
  wire [31:0] _is_aligned_T = io_in_a_bits_address & _GEN_71; // @[Edges.scala 20:16 chipyard.TestHarness.SmallBoomConfig.fir 391138:6]
  wire  is_aligned = _is_aligned_T == 32'h0; // @[Edges.scala 20:24 chipyard.TestHarness.SmallBoomConfig.fir 391139:6]
  wire [1:0] mask_sizeOH_shiftAmount = io_in_a_bits_size[1:0]; // @[OneHot.scala 64:49 chipyard.TestHarness.SmallBoomConfig.fir 391141:6]
  wire [3:0] _mask_sizeOH_T_1 = 4'h1 << mask_sizeOH_shiftAmount; // @[OneHot.scala 65:12 chipyard.TestHarness.SmallBoomConfig.fir 391142:6]
  wire [2:0] mask_sizeOH = _mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81 chipyard.TestHarness.SmallBoomConfig.fir 391144:6]
  wire  _mask_T = io_in_a_bits_size >= 4'h3; // @[Misc.scala 205:21 chipyard.TestHarness.SmallBoomConfig.fir 391145:6]
  wire  mask_size = mask_sizeOH[2]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 391146:6]
  wire  mask_bit = io_in_a_bits_address[2]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 391147:6]
  wire  mask_nbit = ~mask_bit; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 391148:6]
  wire  _mask_acc_T = mask_size & mask_nbit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391150:6]
  wire  mask_acc = _mask_T | _mask_acc_T; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391151:6]
  wire  _mask_acc_T_1 = mask_size & mask_bit; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391153:6]
  wire  mask_acc_1 = _mask_T | _mask_acc_T_1; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391154:6]
  wire  mask_size_1 = mask_sizeOH[1]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 391155:6]
  wire  mask_bit_1 = io_in_a_bits_address[1]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 391156:6]
  wire  mask_nbit_1 = ~mask_bit_1; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 391157:6]
  wire  mask_eq_2 = mask_nbit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391158:6]
  wire  _mask_acc_T_2 = mask_size_1 & mask_eq_2; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391159:6]
  wire  mask_acc_2 = mask_acc | _mask_acc_T_2; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391160:6]
  wire  mask_eq_3 = mask_nbit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391161:6]
  wire  _mask_acc_T_3 = mask_size_1 & mask_eq_3; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391162:6]
  wire  mask_acc_3 = mask_acc | _mask_acc_T_3; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391163:6]
  wire  mask_eq_4 = mask_bit & mask_nbit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391164:6]
  wire  _mask_acc_T_4 = mask_size_1 & mask_eq_4; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391165:6]
  wire  mask_acc_4 = mask_acc_1 | _mask_acc_T_4; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391166:6]
  wire  mask_eq_5 = mask_bit & mask_bit_1; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391167:6]
  wire  _mask_acc_T_5 = mask_size_1 & mask_eq_5; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391168:6]
  wire  mask_acc_5 = mask_acc_1 | _mask_acc_T_5; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391169:6]
  wire  mask_size_2 = mask_sizeOH[0]; // @[Misc.scala 208:26 chipyard.TestHarness.SmallBoomConfig.fir 391170:6]
  wire  mask_bit_2 = io_in_a_bits_address[0]; // @[Misc.scala 209:26 chipyard.TestHarness.SmallBoomConfig.fir 391171:6]
  wire  mask_nbit_2 = ~mask_bit_2; // @[Misc.scala 210:20 chipyard.TestHarness.SmallBoomConfig.fir 391172:6]
  wire  mask_eq_6 = mask_eq_2 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391173:6]
  wire  _mask_acc_T_6 = mask_size_2 & mask_eq_6; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391174:6]
  wire  mask_lo_lo_lo = mask_acc_2 | _mask_acc_T_6; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391175:6]
  wire  mask_eq_7 = mask_eq_2 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391176:6]
  wire  _mask_acc_T_7 = mask_size_2 & mask_eq_7; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391177:6]
  wire  mask_lo_lo_hi = mask_acc_2 | _mask_acc_T_7; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391178:6]
  wire  mask_eq_8 = mask_eq_3 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391179:6]
  wire  _mask_acc_T_8 = mask_size_2 & mask_eq_8; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391180:6]
  wire  mask_lo_hi_lo = mask_acc_3 | _mask_acc_T_8; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391181:6]
  wire  mask_eq_9 = mask_eq_3 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391182:6]
  wire  _mask_acc_T_9 = mask_size_2 & mask_eq_9; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391183:6]
  wire  mask_lo_hi_hi = mask_acc_3 | _mask_acc_T_9; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391184:6]
  wire  mask_eq_10 = mask_eq_4 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391185:6]
  wire  _mask_acc_T_10 = mask_size_2 & mask_eq_10; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391186:6]
  wire  mask_hi_lo_lo = mask_acc_4 | _mask_acc_T_10; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391187:6]
  wire  mask_eq_11 = mask_eq_4 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391188:6]
  wire  _mask_acc_T_11 = mask_size_2 & mask_eq_11; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391189:6]
  wire  mask_hi_lo_hi = mask_acc_4 | _mask_acc_T_11; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391190:6]
  wire  mask_eq_12 = mask_eq_5 & mask_nbit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391191:6]
  wire  _mask_acc_T_12 = mask_size_2 & mask_eq_12; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391192:6]
  wire  mask_hi_hi_lo = mask_acc_5 | _mask_acc_T_12; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391193:6]
  wire  mask_eq_13 = mask_eq_5 & mask_bit_2; // @[Misc.scala 213:27 chipyard.TestHarness.SmallBoomConfig.fir 391194:6]
  wire  _mask_acc_T_13 = mask_size_2 & mask_eq_13; // @[Misc.scala 214:38 chipyard.TestHarness.SmallBoomConfig.fir 391195:6]
  wire  mask_hi_hi_hi = mask_acc_5 | _mask_acc_T_13; // @[Misc.scala 214:29 chipyard.TestHarness.SmallBoomConfig.fir 391196:6]
  wire [7:0] mask = {mask_hi_hi_hi,mask_hi_hi_lo,mask_hi_lo_hi,mask_hi_lo_lo,mask_lo_hi_hi,mask_lo_hi_lo,mask_lo_lo_hi,
    mask_lo_lo_lo}; // @[Cat.scala 30:58 chipyard.TestHarness.SmallBoomConfig.fir 391203:6]
  wire [32:0] _T_7 = {1'b0,$signed(io_in_a_bits_address)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391207:6]
  wire  _T_15 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 81:25 chipyard.TestHarness.SmallBoomConfig.fir 391219:6]
  wire  _T_17 = io_in_a_bits_size <= 4'hc; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 391222:8]
  wire [32:0] _T_26 = $signed(_T_7) & -33'sh101000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391231:8]
  wire  _T_27 = $signed(_T_26) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391232:8]
  wire [31:0] _T_28 = io_in_a_bits_address ^ 32'h3000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391233:8]
  wire [32:0] _T_29 = {1'b0,$signed(_T_28)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391234:8]
  wire [32:0] _T_31 = $signed(_T_29) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391236:8]
  wire  _T_32 = $signed(_T_31) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391237:8]
  wire [31:0] _T_33 = io_in_a_bits_address ^ 32'h10000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391238:8]
  wire [32:0] _T_34 = {1'b0,$signed(_T_33)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391239:8]
  wire [32:0] _T_36 = $signed(_T_34) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391241:8]
  wire  _T_37 = $signed(_T_36) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391242:8]
  wire [31:0] _T_38 = io_in_a_bits_address ^ 32'h2000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391243:8]
  wire [32:0] _T_39 = {1'b0,$signed(_T_38)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391244:8]
  wire [32:0] _T_41 = $signed(_T_39) & -33'sh10000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391246:8]
  wire  _T_42 = $signed(_T_41) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391247:8]
  wire [31:0] _T_43 = io_in_a_bits_address ^ 32'h2010000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391248:8]
  wire [32:0] _T_44 = {1'b0,$signed(_T_43)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391249:8]
  wire [32:0] _T_46 = $signed(_T_44) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391251:8]
  wire  _T_47 = $signed(_T_46) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391252:8]
  wire [31:0] _T_48 = io_in_a_bits_address ^ 32'hc000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391253:8]
  wire [32:0] _T_49 = {1'b0,$signed(_T_48)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391254:8]
  wire [32:0] _T_51 = $signed(_T_49) & -33'sh4000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391256:8]
  wire  _T_52 = $signed(_T_51) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391257:8]
  wire [31:0] _T_53 = io_in_a_bits_address ^ 32'h54000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391258:8]
  wire [32:0] _T_54 = {1'b0,$signed(_T_53)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391259:8]
  wire [32:0] _T_56 = $signed(_T_54) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391261:8]
  wire  _T_57 = $signed(_T_56) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391262:8]
  wire  _T_58 = _T_27 | _T_32; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391263:8]
  wire  _T_65 = 4'h6 == io_in_a_bits_size; // @[Parameters.scala 91:48 chipyard.TestHarness.SmallBoomConfig.fir 391270:8]
  wire [31:0] _T_67 = io_in_a_bits_address ^ 32'h10000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391272:8]
  wire [32:0] _T_68 = {1'b0,$signed(_T_67)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391273:8]
  wire [32:0] _T_70 = $signed(_T_68) & -33'sh1000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391275:8]
  wire  _T_71 = $signed(_T_70) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391276:8]
  wire [31:0] _T_72 = io_in_a_bits_address ^ 32'h80000000; // @[Parameters.scala 137:31 chipyard.TestHarness.SmallBoomConfig.fir 391277:8]
  wire [32:0] _T_73 = {1'b0,$signed(_T_72)}; // @[Parameters.scala 137:49 chipyard.TestHarness.SmallBoomConfig.fir 391278:8]
  wire [32:0] _T_75 = $signed(_T_73) & -33'sh10000000; // @[Parameters.scala 137:52 chipyard.TestHarness.SmallBoomConfig.fir 391280:8]
  wire  _T_76 = $signed(_T_75) == 33'sh0; // @[Parameters.scala 137:67 chipyard.TestHarness.SmallBoomConfig.fir 391281:8]
  wire  _T_77 = _T_71 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391282:8]
  wire  _T_78 = _T_65 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391283:8]
  wire  _T_81 = _T_17 & _T_78; // @[Monitor.scala 82:72 chipyard.TestHarness.SmallBoomConfig.fir 391286:8]
  wire  _T_83 = _T_81 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391288:8]
  wire  _T_84 = ~_T_83; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391289:8]
  wire  _T_147 = ~reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391356:8]
  wire  _T_153 = _mask_T | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391370:8]
  wire  _T_154 = ~_T_153; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391371:8]
  wire  _T_156 = is_aligned | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391377:8]
  wire  _T_157 = ~_T_156; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391378:8]
  wire [7:0] _T_162 = ~io_in_a_bits_mask; // @[Monitor.scala 88:18 chipyard.TestHarness.SmallBoomConfig.fir 391391:8]
  wire  _T_163 = _T_162 == 8'h0; // @[Monitor.scala 88:31 chipyard.TestHarness.SmallBoomConfig.fir 391392:8]
  wire  _T_165 = _T_163 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391394:8]
  wire  _T_166 = ~_T_165; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391395:8]
  wire  _T_171 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 92:25 chipyard.TestHarness.SmallBoomConfig.fir 391409:6]
  wire  _T_331 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 104:25 chipyard.TestHarness.SmallBoomConfig.fir 391607:6]
  wire  _T_339 = _T_17 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391616:8]
  wire  _T_340 = ~_T_339; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391617:8]
  wire  _T_350 = _T_17 & _T_32; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391631:8]
  wire  _T_352 = io_in_a_bits_size <= 4'h6; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 391633:8]
  wire  _T_395 = _T_27 | _T_37; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391676:8]
  wire  _T_396 = _T_395 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391677:8]
  wire  _T_397 = _T_396 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391678:8]
  wire  _T_398 = _T_397 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391679:8]
  wire  _T_399 = _T_398 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391680:8]
  wire  _T_400 = _T_399 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391681:8]
  wire  _T_401 = _T_400 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391682:8]
  wire  _T_402 = _T_352 & _T_401; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391683:8]
  wire  _T_404 = _T_350 | _T_402; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 391685:8]
  wire  _T_406 = _T_404 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391687:8]
  wire  _T_407 = ~_T_406; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391688:8]
  wire  _T_418 = io_in_a_bits_mask == mask; // @[Monitor.scala 110:30 chipyard.TestHarness.SmallBoomConfig.fir 391715:8]
  wire  _T_420 = _T_418 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391717:8]
  wire  _T_421 = ~_T_420; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391718:8]
  wire  _T_426 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 114:25 chipyard.TestHarness.SmallBoomConfig.fir 391732:6]
  wire  _T_482 = _T_27 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391789:8]
  wire  _T_483 = _T_482 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391790:8]
  wire  _T_484 = _T_483 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391791:8]
  wire  _T_485 = _T_484 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391792:8]
  wire  _T_486 = _T_485 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391793:8]
  wire  _T_487 = _T_486 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 391794:8]
  wire  _T_488 = _T_352 & _T_487; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 391795:8]
  wire  _T_497 = _T_350 | _T_488; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 391804:8]
  wire  _T_499 = _T_17 & _T_497; // @[Monitor.scala 115:71 chipyard.TestHarness.SmallBoomConfig.fir 391806:8]
  wire  _T_501 = _T_499 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391808:8]
  wire  _T_502 = ~_T_501; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391809:8]
  wire  _T_517 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 122:25 chipyard.TestHarness.SmallBoomConfig.fir 391845:6]
  wire [7:0] _T_604 = ~mask; // @[Monitor.scala 127:33 chipyard.TestHarness.SmallBoomConfig.fir 391949:8]
  wire [7:0] _T_605 = io_in_a_bits_mask & _T_604; // @[Monitor.scala 127:31 chipyard.TestHarness.SmallBoomConfig.fir 391950:8]
  wire  _T_606 = _T_605 == 8'h0; // @[Monitor.scala 127:40 chipyard.TestHarness.SmallBoomConfig.fir 391951:8]
  wire  _T_608 = _T_606 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391953:8]
  wire  _T_609 = ~_T_608; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391954:8]
  wire  _T_610 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 130:25 chipyard.TestHarness.SmallBoomConfig.fir 391960:6]
  wire  _T_618 = io_in_a_bits_size <= 4'h3; // @[Parameters.scala 92:42 chipyard.TestHarness.SmallBoomConfig.fir 391969:8]
  wire  _T_662 = _T_58 | _T_42; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392013:8]
  wire  _T_663 = _T_662 | _T_47; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392014:8]
  wire  _T_664 = _T_663 | _T_52; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392015:8]
  wire  _T_665 = _T_664 | _T_71; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392016:8]
  wire  _T_666 = _T_665 | _T_57; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392017:8]
  wire  _T_667 = _T_666 | _T_76; // @[Parameters.scala 671:42 chipyard.TestHarness.SmallBoomConfig.fir 392018:8]
  wire  _T_668 = _T_618 & _T_667; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 392019:8]
  wire  _T_678 = _T_17 & _T_668; // @[Monitor.scala 131:74 chipyard.TestHarness.SmallBoomConfig.fir 392029:8]
  wire  _T_680 = _T_678 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392031:8]
  wire  _T_681 = ~_T_680; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392032:8]
  wire  _T_696 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 138:25 chipyard.TestHarness.SmallBoomConfig.fir 392068:6]
  wire  _T_782 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 146:25 chipyard.TestHarness.SmallBoomConfig.fir 392176:6]
  wire  _T_851 = _T_352 & _T_77; // @[Parameters.scala 670:56 chipyard.TestHarness.SmallBoomConfig.fir 392246:8]
  wire  _T_854 = _T_350 | _T_851; // @[Parameters.scala 672:30 chipyard.TestHarness.SmallBoomConfig.fir 392249:8]
  wire  _T_855 = _T_17 & _T_854; // @[Monitor.scala 147:68 chipyard.TestHarness.SmallBoomConfig.fir 392250:8]
  wire  _T_857 = _T_855 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392252:8]
  wire  _T_858 = ~_T_857; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392253:8]
  wire  _T_877 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 42:24 chipyard.TestHarness.SmallBoomConfig.fir 392299:6]
  wire  _T_879 = _T_877 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392301:6]
  wire  _T_880 = ~_T_879; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392302:6]
  wire  _source_ok_T_1 = ~io_in_d_bits_source; // @[Parameters.scala 46:9 chipyard.TestHarness.SmallBoomConfig.fir 392307:6]
  wire  _T_881 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 310:25 chipyard.TestHarness.SmallBoomConfig.fir 392312:6]
  wire  _T_883 = _source_ok_T_1 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392315:8]
  wire  _T_884 = ~_T_883; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392316:8]
  wire  _T_885 = io_in_d_bits_size >= 4'h3; // @[Monitor.scala 312:27 chipyard.TestHarness.SmallBoomConfig.fir 392321:8]
  wire  _T_887 = _T_885 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392323:8]
  wire  _T_888 = ~_T_887; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392324:8]
  wire  _T_889 = io_in_d_bits_param == 2'h0; // @[Monitor.scala 313:28 chipyard.TestHarness.SmallBoomConfig.fir 392329:8]
  wire  _T_891 = _T_889 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392331:8]
  wire  _T_892 = ~_T_891; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392332:8]
  wire  _T_893 = ~io_in_d_bits_corrupt; // @[Monitor.scala 314:15 chipyard.TestHarness.SmallBoomConfig.fir 392337:8]
  wire  _T_895 = _T_893 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392339:8]
  wire  _T_896 = ~_T_895; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392340:8]
  wire  _T_897 = ~io_in_d_bits_denied; // @[Monitor.scala 315:15 chipyard.TestHarness.SmallBoomConfig.fir 392345:8]
  wire  _T_899 = _T_897 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392347:8]
  wire  _T_900 = ~_T_899; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392348:8]
  wire  _T_901 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 318:25 chipyard.TestHarness.SmallBoomConfig.fir 392354:6]
  wire  _T_912 = io_in_d_bits_param <= 2'h2; // @[Bundles.scala 102:26 chipyard.TestHarness.SmallBoomConfig.fir 392378:8]
  wire  _T_914 = _T_912 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392380:8]
  wire  _T_915 = ~_T_914; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392381:8]
  wire  _T_916 = io_in_d_bits_param != 2'h2; // @[Monitor.scala 323:28 chipyard.TestHarness.SmallBoomConfig.fir 392386:8]
  wire  _T_918 = _T_916 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392388:8]
  wire  _T_919 = ~_T_918; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392389:8]
  wire  _T_929 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 328:25 chipyard.TestHarness.SmallBoomConfig.fir 392412:6]
  wire  _T_949 = _T_897 | io_in_d_bits_corrupt; // @[Monitor.scala 334:30 chipyard.TestHarness.SmallBoomConfig.fir 392453:8]
  wire  _T_951 = _T_949 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392455:8]
  wire  _T_952 = ~_T_951; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392456:8]
  wire  _T_958 = io_in_d_bits_opcode == 3'h0; // @[Monitor.scala 338:25 chipyard.TestHarness.SmallBoomConfig.fir 392471:6]
  wire  _T_975 = io_in_d_bits_opcode == 3'h1; // @[Monitor.scala 346:25 chipyard.TestHarness.SmallBoomConfig.fir 392506:6]
  wire  _T_993 = io_in_d_bits_opcode == 3'h2; // @[Monitor.scala 354:25 chipyard.TestHarness.SmallBoomConfig.fir 392542:6]
  wire  _a_first_T = io_in_a_ready & io_in_a_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 392608:4]
  wire [8:0] a_first_beats1_decode = is_aligned_mask[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 392613:4]
  wire  a_first_beats1_opdata = ~io_in_a_bits_opcode[2]; // @[Edges.scala 91:28 chipyard.TestHarness.SmallBoomConfig.fir 392615:4]
  reg [8:0] a_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392617:4]
  wire [8:0] a_first_counter1 = a_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392619:4]
  wire  a_first = a_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392620:4]
  reg [2:0] opcode; // @[Monitor.scala 384:22 chipyard.TestHarness.SmallBoomConfig.fir 392631:4]
  reg [3:0] size; // @[Monitor.scala 386:22 chipyard.TestHarness.SmallBoomConfig.fir 392633:4]
  reg [31:0] address; // @[Monitor.scala 388:22 chipyard.TestHarness.SmallBoomConfig.fir 392635:4]
  wire  _T_1022 = ~a_first; // @[Monitor.scala 389:22 chipyard.TestHarness.SmallBoomConfig.fir 392636:4]
  wire  _T_1023 = io_in_a_valid & _T_1022; // @[Monitor.scala 389:19 chipyard.TestHarness.SmallBoomConfig.fir 392637:4]
  wire  _T_1024 = io_in_a_bits_opcode == opcode; // @[Monitor.scala 390:32 chipyard.TestHarness.SmallBoomConfig.fir 392639:6]
  wire  _T_1026 = _T_1024 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392641:6]
  wire  _T_1027 = ~_T_1026; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392642:6]
  wire  _T_1032 = io_in_a_bits_size == size; // @[Monitor.scala 392:32 chipyard.TestHarness.SmallBoomConfig.fir 392655:6]
  wire  _T_1034 = _T_1032 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392657:6]
  wire  _T_1035 = ~_T_1034; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392658:6]
  wire  _T_1040 = io_in_a_bits_address == address; // @[Monitor.scala 394:32 chipyard.TestHarness.SmallBoomConfig.fir 392671:6]
  wire  _T_1042 = _T_1040 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392673:6]
  wire  _T_1043 = ~_T_1042; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392674:6]
  wire  _T_1045 = _a_first_T & a_first; // @[Monitor.scala 396:20 chipyard.TestHarness.SmallBoomConfig.fir 392681:4]
  wire  _d_first_T = io_in_d_ready & io_in_d_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 392689:4]
  wire [26:0] _d_first_beats1_decode_T_1 = 27'hfff << io_in_d_bits_size; // @[package.scala 234:77 chipyard.TestHarness.SmallBoomConfig.fir 392691:4]
  wire [11:0] _d_first_beats1_decode_T_3 = ~_d_first_beats1_decode_T_1[11:0]; // @[package.scala 234:46 chipyard.TestHarness.SmallBoomConfig.fir 392693:4]
  wire [8:0] d_first_beats1_decode = _d_first_beats1_decode_T_3[11:3]; // @[Edges.scala 219:59 chipyard.TestHarness.SmallBoomConfig.fir 392694:4]
  wire  d_first_beats1_opdata = io_in_d_bits_opcode[0]; // @[Edges.scala 105:36 chipyard.TestHarness.SmallBoomConfig.fir 392695:4]
  reg [8:0] d_first_counter; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392697:4]
  wire [8:0] d_first_counter1 = d_first_counter - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392699:4]
  wire  d_first = d_first_counter == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392700:4]
  reg [2:0] opcode_1; // @[Monitor.scala 535:22 chipyard.TestHarness.SmallBoomConfig.fir 392711:4]
  reg [1:0] param_1; // @[Monitor.scala 536:22 chipyard.TestHarness.SmallBoomConfig.fir 392712:4]
  reg [3:0] size_1; // @[Monitor.scala 537:22 chipyard.TestHarness.SmallBoomConfig.fir 392713:4]
  reg  source_1; // @[Monitor.scala 538:22 chipyard.TestHarness.SmallBoomConfig.fir 392714:4]
  reg [2:0] sink; // @[Monitor.scala 539:22 chipyard.TestHarness.SmallBoomConfig.fir 392715:4]
  reg  denied; // @[Monitor.scala 540:22 chipyard.TestHarness.SmallBoomConfig.fir 392716:4]
  wire  _T_1046 = ~d_first; // @[Monitor.scala 541:22 chipyard.TestHarness.SmallBoomConfig.fir 392717:4]
  wire  _T_1047 = io_in_d_valid & _T_1046; // @[Monitor.scala 541:19 chipyard.TestHarness.SmallBoomConfig.fir 392718:4]
  wire  _T_1048 = io_in_d_bits_opcode == opcode_1; // @[Monitor.scala 542:29 chipyard.TestHarness.SmallBoomConfig.fir 392720:6]
  wire  _T_1050 = _T_1048 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392722:6]
  wire  _T_1051 = ~_T_1050; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392723:6]
  wire  _T_1052 = io_in_d_bits_param == param_1; // @[Monitor.scala 543:29 chipyard.TestHarness.SmallBoomConfig.fir 392728:6]
  wire  _T_1054 = _T_1052 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392730:6]
  wire  _T_1055 = ~_T_1054; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392731:6]
  wire  _T_1056 = io_in_d_bits_size == size_1; // @[Monitor.scala 544:29 chipyard.TestHarness.SmallBoomConfig.fir 392736:6]
  wire  _T_1058 = _T_1056 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392738:6]
  wire  _T_1059 = ~_T_1058; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392739:6]
  wire  _T_1060 = io_in_d_bits_source == source_1; // @[Monitor.scala 545:29 chipyard.TestHarness.SmallBoomConfig.fir 392744:6]
  wire  _T_1062 = _T_1060 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392746:6]
  wire  _T_1063 = ~_T_1062; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392747:6]
  wire  _T_1064 = io_in_d_bits_sink == sink; // @[Monitor.scala 546:29 chipyard.TestHarness.SmallBoomConfig.fir 392752:6]
  wire  _T_1066 = _T_1064 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392754:6]
  wire  _T_1067 = ~_T_1066; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392755:6]
  wire  _T_1068 = io_in_d_bits_denied == denied; // @[Monitor.scala 547:29 chipyard.TestHarness.SmallBoomConfig.fir 392760:6]
  wire  _T_1070 = _T_1068 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392762:6]
  wire  _T_1071 = ~_T_1070; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392763:6]
  wire  _T_1073 = _d_first_T & d_first; // @[Monitor.scala 549:20 chipyard.TestHarness.SmallBoomConfig.fir 392770:4]
  reg  inflight; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 392779:4]
  reg [3:0] inflight_opcodes; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 392780:4]
  reg [7:0] inflight_sizes; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 392781:4]
  reg [8:0] a_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392791:4]
  wire [8:0] a_first_counter1_1 = a_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392793:4]
  wire  a_first_1 = a_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392794:4]
  reg [8:0] d_first_counter_1; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392813:4]
  wire [8:0] d_first_counter1_1 = d_first_counter_1 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 392815:4]
  wire  d_first_1 = d_first_counter_1 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 392816:4]
  wire [2:0] _GEN_72 = {io_in_d_bits_source, 2'h0}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 392837:4]
  wire [3:0] _a_opcode_lookup_T = {{1'd0}, _GEN_72}; // @[Monitor.scala 634:69 chipyard.TestHarness.SmallBoomConfig.fir 392837:4]
  wire [3:0] _a_opcode_lookup_T_1 = inflight_opcodes >> _a_opcode_lookup_T; // @[Monitor.scala 634:44 chipyard.TestHarness.SmallBoomConfig.fir 392838:4]
  wire [15:0] _a_opcode_lookup_T_5 = 16'h10 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 392842:4]
  wire [15:0] _GEN_73 = {{12'd0}, _a_opcode_lookup_T_1}; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 392843:4]
  wire [15:0] _a_opcode_lookup_T_6 = _GEN_73 & _a_opcode_lookup_T_5; // @[Monitor.scala 634:97 chipyard.TestHarness.SmallBoomConfig.fir 392843:4]
  wire [15:0] _a_opcode_lookup_T_7 = {{1'd0}, _a_opcode_lookup_T_6[15:1]}; // @[Monitor.scala 634:152 chipyard.TestHarness.SmallBoomConfig.fir 392844:4]
  wire [3:0] _a_size_lookup_T = {io_in_d_bits_source, 3'h0}; // @[Monitor.scala 638:65 chipyard.TestHarness.SmallBoomConfig.fir 392848:4]
  wire [7:0] _a_size_lookup_T_1 = inflight_sizes >> _a_size_lookup_T; // @[Monitor.scala 638:40 chipyard.TestHarness.SmallBoomConfig.fir 392849:4]
  wire [15:0] _a_size_lookup_T_5 = 16'h100 - 16'h1; // @[Monitor.scala 609:57 chipyard.TestHarness.SmallBoomConfig.fir 392853:4]
  wire [15:0] _GEN_75 = {{8'd0}, _a_size_lookup_T_1}; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 392854:4]
  wire [15:0] _a_size_lookup_T_6 = _GEN_75 & _a_size_lookup_T_5; // @[Monitor.scala 638:91 chipyard.TestHarness.SmallBoomConfig.fir 392854:4]
  wire [15:0] _a_size_lookup_T_7 = {{1'd0}, _a_size_lookup_T_6[15:1]}; // @[Monitor.scala 638:144 chipyard.TestHarness.SmallBoomConfig.fir 392855:4]
  wire  _T_1074 = io_in_a_valid & a_first_1; // @[Monitor.scala 648:26 chipyard.TestHarness.SmallBoomConfig.fir 392879:4]
  wire [1:0] _GEN_15 = _T_1074 ? 2'h1 : 2'h0; // @[Monitor.scala 648:71 chipyard.TestHarness.SmallBoomConfig.fir 392881:4 Monitor.scala 649:22 chipyard.TestHarness.SmallBoomConfig.fir 392883:6 chipyard.TestHarness.SmallBoomConfig.fir 392830:4]
  wire  _T_1077 = _a_first_T & a_first_1; // @[Monitor.scala 652:27 chipyard.TestHarness.SmallBoomConfig.fir 392886:4]
  wire [3:0] _a_opcodes_set_interm_T = {io_in_a_bits_opcode, 1'h0}; // @[Monitor.scala 654:53 chipyard.TestHarness.SmallBoomConfig.fir 392891:6]
  wire [3:0] _a_opcodes_set_interm_T_1 = _a_opcodes_set_interm_T | 4'h1; // @[Monitor.scala 654:61 chipyard.TestHarness.SmallBoomConfig.fir 392892:6]
  wire [4:0] _a_sizes_set_interm_T = {io_in_a_bits_size, 1'h0}; // @[Monitor.scala 655:51 chipyard.TestHarness.SmallBoomConfig.fir 392894:6]
  wire [4:0] _a_sizes_set_interm_T_1 = _a_sizes_set_interm_T | 5'h1; // @[Monitor.scala 655:59 chipyard.TestHarness.SmallBoomConfig.fir 392895:6]
  wire [3:0] a_opcodes_set_interm = _T_1077 ? _a_opcodes_set_interm_T_1 : 4'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392888:4 Monitor.scala 654:28 chipyard.TestHarness.SmallBoomConfig.fir 392893:6 chipyard.TestHarness.SmallBoomConfig.fir 392876:4]
  wire [18:0] _a_opcodes_set_T_1 = {{15'd0}, a_opcodes_set_interm}; // @[Monitor.scala 656:54 chipyard.TestHarness.SmallBoomConfig.fir 392898:6]
  wire [4:0] a_sizes_set_interm = _T_1077 ? _a_sizes_set_interm_T_1 : 5'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392888:4 Monitor.scala 655:28 chipyard.TestHarness.SmallBoomConfig.fir 392896:6 chipyard.TestHarness.SmallBoomConfig.fir 392878:4]
  wire [19:0] _a_sizes_set_T_1 = {{15'd0}, a_sizes_set_interm}; // @[Monitor.scala 657:52 chipyard.TestHarness.SmallBoomConfig.fir 392901:6]
  wire  _T_1081 = ~inflight; // @[Monitor.scala 658:17 chipyard.TestHarness.SmallBoomConfig.fir 392905:6]
  wire  _T_1083 = _T_1081 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392907:6]
  wire  _T_1084 = ~_T_1083; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392908:6]
  wire [1:0] _GEN_16 = _T_1077 ? 2'h1 : 2'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392888:4 Monitor.scala 653:28 chipyard.TestHarness.SmallBoomConfig.fir 392890:6 chipyard.TestHarness.SmallBoomConfig.fir 392828:4]
  wire [18:0] _GEN_19 = _T_1077 ? _a_opcodes_set_T_1 : 19'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392888:4 Monitor.scala 656:28 chipyard.TestHarness.SmallBoomConfig.fir 392899:6 chipyard.TestHarness.SmallBoomConfig.fir 392832:4]
  wire [19:0] _GEN_20 = _T_1077 ? _a_sizes_set_T_1 : 20'h0; // @[Monitor.scala 652:72 chipyard.TestHarness.SmallBoomConfig.fir 392888:4 Monitor.scala 657:28 chipyard.TestHarness.SmallBoomConfig.fir 392902:6 chipyard.TestHarness.SmallBoomConfig.fir 392834:4]
  wire  _T_1085 = io_in_d_valid & d_first_1; // @[Monitor.scala 671:26 chipyard.TestHarness.SmallBoomConfig.fir 392923:4]
  wire  _T_1087 = ~_T_881; // @[Monitor.scala 671:74 chipyard.TestHarness.SmallBoomConfig.fir 392925:4]
  wire  _T_1088 = _T_1085 & _T_1087; // @[Monitor.scala 671:71 chipyard.TestHarness.SmallBoomConfig.fir 392926:4]
  wire [1:0] _d_clr_wo_ready_T = 2'h1 << io_in_d_bits_source; // @[OneHot.scala 58:35 chipyard.TestHarness.SmallBoomConfig.fir 392928:6]
  wire [1:0] _GEN_21 = _T_1088 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 671:90 chipyard.TestHarness.SmallBoomConfig.fir 392927:4 Monitor.scala 672:22 chipyard.TestHarness.SmallBoomConfig.fir 392929:6 chipyard.TestHarness.SmallBoomConfig.fir 392917:4]
  wire  _T_1090 = _d_first_T & d_first_1; // @[Monitor.scala 675:27 chipyard.TestHarness.SmallBoomConfig.fir 392932:4]
  wire  _T_1093 = _T_1090 & _T_1087; // @[Monitor.scala 675:72 chipyard.TestHarness.SmallBoomConfig.fir 392935:4]
  wire [30:0] _GEN_78 = {{15'd0}, _a_opcode_lookup_T_5}; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 392944:6]
  wire [30:0] _d_opcodes_clr_T_5 = _GEN_78 << _a_opcode_lookup_T; // @[Monitor.scala 677:76 chipyard.TestHarness.SmallBoomConfig.fir 392944:6]
  wire [30:0] _GEN_79 = {{15'd0}, _a_size_lookup_T_5}; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 392951:6]
  wire [30:0] _d_sizes_clr_T_5 = _GEN_79 << _a_size_lookup_T; // @[Monitor.scala 678:74 chipyard.TestHarness.SmallBoomConfig.fir 392951:6]
  wire [1:0] _GEN_22 = _T_1093 ? _d_clr_wo_ready_T : 2'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 392936:4 Monitor.scala 676:21 chipyard.TestHarness.SmallBoomConfig.fir 392938:6 chipyard.TestHarness.SmallBoomConfig.fir 392915:4]
  wire [30:0] _GEN_23 = _T_1093 ? _d_opcodes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 392936:4 Monitor.scala 677:21 chipyard.TestHarness.SmallBoomConfig.fir 392945:6 chipyard.TestHarness.SmallBoomConfig.fir 392919:4]
  wire [30:0] _GEN_24 = _T_1093 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 675:91 chipyard.TestHarness.SmallBoomConfig.fir 392936:4 Monitor.scala 678:21 chipyard.TestHarness.SmallBoomConfig.fir 392952:6 chipyard.TestHarness.SmallBoomConfig.fir 392921:4]
  wire  same_cycle_resp = _T_1074 & _source_ok_T_1; // @[Monitor.scala 681:88 chipyard.TestHarness.SmallBoomConfig.fir 392962:6]
  wire  _T_1098 = inflight >> io_in_d_bits_source; // @[Monitor.scala 682:25 chipyard.TestHarness.SmallBoomConfig.fir 392963:6]
  wire  _T_1100 = _T_1098 | same_cycle_resp; // @[Monitor.scala 682:49 chipyard.TestHarness.SmallBoomConfig.fir 392965:6]
  wire  _T_1102 = _T_1100 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392967:6]
  wire  _T_1103 = ~_T_1102; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392968:6]
  wire [2:0] _GEN_27 = 3'h2 == io_in_a_bits_opcode ? 3'h1 : 3'h0; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8]
  wire [2:0] _GEN_28 = 3'h3 == io_in_a_bits_opcode ? 3'h1 : _GEN_27; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8]
  wire [2:0] _GEN_29 = 3'h4 == io_in_a_bits_opcode ? 3'h1 : _GEN_28; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8]
  wire [2:0] _GEN_30 = 3'h5 == io_in_a_bits_opcode ? 3'h2 : _GEN_29; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8]
  wire [2:0] _GEN_31 = 3'h6 == io_in_a_bits_opcode ? 3'h4 : _GEN_30; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8]
  wire [2:0] _GEN_32 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_31; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8 Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8]
  wire  _T_1104 = io_in_d_bits_opcode == _GEN_32; // @[Monitor.scala 685:38 chipyard.TestHarness.SmallBoomConfig.fir 392974:8]
  wire [2:0] _GEN_39 = 3'h6 == io_in_a_bits_opcode ? 3'h5 : _GEN_30; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 392975:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 392975:8]
  wire [2:0] _GEN_40 = 3'h7 == io_in_a_bits_opcode ? 3'h4 : _GEN_39; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 392975:8 Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 392975:8]
  wire  _T_1105 = io_in_d_bits_opcode == _GEN_40; // @[Monitor.scala 686:39 chipyard.TestHarness.SmallBoomConfig.fir 392975:8]
  wire  _T_1106 = _T_1104 | _T_1105; // @[Monitor.scala 685:77 chipyard.TestHarness.SmallBoomConfig.fir 392976:8]
  wire  _T_1108 = _T_1106 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392978:8]
  wire  _T_1109 = ~_T_1108; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392979:8]
  wire  _T_1110 = io_in_a_bits_size == io_in_d_bits_size; // @[Monitor.scala 687:36 chipyard.TestHarness.SmallBoomConfig.fir 392984:8]
  wire  _T_1112 = _T_1110 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392986:8]
  wire  _T_1113 = ~_T_1112; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392987:8]
  wire [3:0] a_opcode_lookup = _a_opcode_lookup_T_7[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392835:4 Monitor.scala 634:21 chipyard.TestHarness.SmallBoomConfig.fir 392845:4]
  wire [2:0] _GEN_43 = 3'h2 == a_opcode_lookup[2:0] ? 3'h1 : 3'h0; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8]
  wire [2:0] _GEN_44 = 3'h3 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_43; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8]
  wire [2:0] _GEN_45 = 3'h4 == a_opcode_lookup[2:0] ? 3'h1 : _GEN_44; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8]
  wire [2:0] _GEN_46 = 3'h5 == a_opcode_lookup[2:0] ? 3'h2 : _GEN_45; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8]
  wire [2:0] _GEN_47 = 3'h6 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_46; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8]
  wire [2:0] _GEN_48 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_47; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8 Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8]
  wire  _T_1115 = io_in_d_bits_opcode == _GEN_48; // @[Monitor.scala 689:38 chipyard.TestHarness.SmallBoomConfig.fir 392995:8]
  wire [2:0] _GEN_55 = 3'h6 == a_opcode_lookup[2:0] ? 3'h5 : _GEN_46; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 392997:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 392997:8]
  wire [2:0] _GEN_56 = 3'h7 == a_opcode_lookup[2:0] ? 3'h4 : _GEN_55; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 392997:8 Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 392997:8]
  wire  _T_1117 = io_in_d_bits_opcode == _GEN_56; // @[Monitor.scala 690:38 chipyard.TestHarness.SmallBoomConfig.fir 392997:8]
  wire  _T_1118 = _T_1115 | _T_1117; // @[Monitor.scala 689:72 chipyard.TestHarness.SmallBoomConfig.fir 392998:8]
  wire  _T_1120 = _T_1118 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393000:8]
  wire  _T_1121 = ~_T_1120; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393001:8]
  wire [7:0] a_size_lookup = _a_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392846:4 Monitor.scala 638:19 chipyard.TestHarness.SmallBoomConfig.fir 392856:4]
  wire [7:0] _GEN_80 = {{4'd0}, io_in_d_bits_size}; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 393006:8]
  wire  _T_1122 = _GEN_80 == a_size_lookup; // @[Monitor.scala 691:36 chipyard.TestHarness.SmallBoomConfig.fir 393006:8]
  wire  _T_1124 = _T_1122 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393008:8]
  wire  _T_1125 = ~_T_1124; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393009:8]
  wire  _T_1127 = _T_1085 & a_first_1; // @[Monitor.scala 694:36 chipyard.TestHarness.SmallBoomConfig.fir 393017:4]
  wire  _T_1128 = _T_1127 & io_in_a_valid; // @[Monitor.scala 694:47 chipyard.TestHarness.SmallBoomConfig.fir 393018:4]
  wire  _T_1130 = _T_1128 & _source_ok_T_1; // @[Monitor.scala 694:65 chipyard.TestHarness.SmallBoomConfig.fir 393020:4]
  wire  _T_1132 = _T_1130 & _T_1087; // @[Monitor.scala 694:116 chipyard.TestHarness.SmallBoomConfig.fir 393022:4]
  wire  _T_1133 = ~io_in_d_ready; // @[Monitor.scala 695:15 chipyard.TestHarness.SmallBoomConfig.fir 393024:6]
  wire  _T_1134 = _T_1133 | io_in_a_ready; // @[Monitor.scala 695:32 chipyard.TestHarness.SmallBoomConfig.fir 393025:6]
  wire  _T_1136 = _T_1134 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393027:6]
  wire  _T_1137 = ~_T_1136; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393028:6]
  wire  a_set_wo_ready = _GEN_15[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392829:4]
  wire  d_clr_wo_ready = _GEN_21[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392916:4]
  wire  _T_1138 = a_set_wo_ready != d_clr_wo_ready; // @[Monitor.scala 699:29 chipyard.TestHarness.SmallBoomConfig.fir 393034:4]
  wire  _T_1139 = |a_set_wo_ready; // @[Monitor.scala 699:67 chipyard.TestHarness.SmallBoomConfig.fir 393035:4]
  wire  _T_1140 = ~_T_1139; // @[Monitor.scala 699:51 chipyard.TestHarness.SmallBoomConfig.fir 393036:4]
  wire  _T_1141 = _T_1138 | _T_1140; // @[Monitor.scala 699:48 chipyard.TestHarness.SmallBoomConfig.fir 393037:4]
  wire  _T_1143 = _T_1141 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393039:4]
  wire  _T_1144 = ~_T_1143; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393040:4]
  wire  a_set = _GEN_16[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392827:4]
  wire  _inflight_T = inflight | a_set; // @[Monitor.scala 702:27 chipyard.TestHarness.SmallBoomConfig.fir 393045:4]
  wire  d_clr = _GEN_22[0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392914:4]
  wire  _inflight_T_1 = ~d_clr; // @[Monitor.scala 702:38 chipyard.TestHarness.SmallBoomConfig.fir 393046:4]
  wire  _inflight_T_2 = _inflight_T & _inflight_T_1; // @[Monitor.scala 702:36 chipyard.TestHarness.SmallBoomConfig.fir 393047:4]
  wire [3:0] a_opcodes_set = _GEN_19[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392831:4]
  wire [3:0] _inflight_opcodes_T = inflight_opcodes | a_opcodes_set; // @[Monitor.scala 703:43 chipyard.TestHarness.SmallBoomConfig.fir 393049:4]
  wire [3:0] d_opcodes_clr = _GEN_23[3:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392918:4]
  wire [3:0] _inflight_opcodes_T_1 = ~d_opcodes_clr; // @[Monitor.scala 703:62 chipyard.TestHarness.SmallBoomConfig.fir 393050:4]
  wire [3:0] _inflight_opcodes_T_2 = _inflight_opcodes_T & _inflight_opcodes_T_1; // @[Monitor.scala 703:60 chipyard.TestHarness.SmallBoomConfig.fir 393051:4]
  wire [7:0] a_sizes_set = _GEN_20[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392833:4]
  wire [7:0] _inflight_sizes_T = inflight_sizes | a_sizes_set; // @[Monitor.scala 704:39 chipyard.TestHarness.SmallBoomConfig.fir 393053:4]
  wire [7:0] d_sizes_clr = _GEN_24[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 392920:4]
  wire [7:0] _inflight_sizes_T_1 = ~d_sizes_clr; // @[Monitor.scala 704:56 chipyard.TestHarness.SmallBoomConfig.fir 393054:4]
  wire [7:0] _inflight_sizes_T_2 = _inflight_sizes_T & _inflight_sizes_T_1; // @[Monitor.scala 704:54 chipyard.TestHarness.SmallBoomConfig.fir 393055:4]
  reg [31:0] watchdog; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 393057:4]
  wire  _T_1145 = |inflight; // @[Monitor.scala 709:26 chipyard.TestHarness.SmallBoomConfig.fir 393060:4]
  wire  _T_1146 = ~_T_1145; // @[Monitor.scala 709:16 chipyard.TestHarness.SmallBoomConfig.fir 393061:4]
  wire  _T_1147 = plusarg_reader_out == 32'h0; // @[Monitor.scala 709:39 chipyard.TestHarness.SmallBoomConfig.fir 393062:4]
  wire  _T_1148 = _T_1146 | _T_1147; // @[Monitor.scala 709:30 chipyard.TestHarness.SmallBoomConfig.fir 393063:4]
  wire  _T_1149 = watchdog < plusarg_reader_out; // @[Monitor.scala 709:59 chipyard.TestHarness.SmallBoomConfig.fir 393064:4]
  wire  _T_1150 = _T_1148 | _T_1149; // @[Monitor.scala 709:47 chipyard.TestHarness.SmallBoomConfig.fir 393065:4]
  wire  _T_1152 = _T_1150 | reset; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393067:4]
  wire  _T_1153 = ~_T_1152; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393068:4]
  wire [31:0] _watchdog_T_1 = watchdog + 32'h1; // @[Monitor.scala 711:26 chipyard.TestHarness.SmallBoomConfig.fir 393074:4]
  wire  _T_1156 = _a_first_T | _d_first_T; // @[Monitor.scala 712:27 chipyard.TestHarness.SmallBoomConfig.fir 393078:4]
  reg [7:0] inflight_sizes_1; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 393084:4]
  reg [8:0] d_first_counter_2; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 393119:4]
  wire [8:0] d_first_counter1_2 = d_first_counter_2 - 9'h1; // @[Edges.scala 229:28 chipyard.TestHarness.SmallBoomConfig.fir 393121:4]
  wire  d_first_2 = d_first_counter_2 == 9'h0; // @[Edges.scala 230:25 chipyard.TestHarness.SmallBoomConfig.fir 393122:4]
  wire [7:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _a_size_lookup_T; // @[Monitor.scala 747:42 chipyard.TestHarness.SmallBoomConfig.fir 393155:4]
  wire [15:0] _GEN_84 = {{8'd0}, _c_size_lookup_T_1}; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 393160:4]
  wire [15:0] _c_size_lookup_T_6 = _GEN_84 & _a_size_lookup_T_5; // @[Monitor.scala 747:93 chipyard.TestHarness.SmallBoomConfig.fir 393160:4]
  wire [15:0] _c_size_lookup_T_7 = {{1'd0}, _c_size_lookup_T_6[15:1]}; // @[Monitor.scala 747:146 chipyard.TestHarness.SmallBoomConfig.fir 393161:4]
  wire  _T_1174 = io_in_d_valid & d_first_2; // @[Monitor.scala 779:26 chipyard.TestHarness.SmallBoomConfig.fir 393239:4]
  wire  _T_1176 = _T_1174 & _T_881; // @[Monitor.scala 779:71 chipyard.TestHarness.SmallBoomConfig.fir 393241:4]
  wire  _T_1178 = _d_first_T & d_first_2; // @[Monitor.scala 783:27 chipyard.TestHarness.SmallBoomConfig.fir 393247:4]
  wire  _T_1180 = _T_1178 & _T_881; // @[Monitor.scala 783:72 chipyard.TestHarness.SmallBoomConfig.fir 393249:4]
  wire [30:0] _GEN_69 = _T_1180 ? _d_sizes_clr_T_5 : 31'h0; // @[Monitor.scala 783:90 chipyard.TestHarness.SmallBoomConfig.fir 393250:4 Monitor.scala 786:21 chipyard.TestHarness.SmallBoomConfig.fir 393266:6 chipyard.TestHarness.SmallBoomConfig.fir 393237:4]
  wire  _T_1184 = 1'h0 >> io_in_d_bits_source; // @[Monitor.scala 791:25 chipyard.TestHarness.SmallBoomConfig.fir 393285:6]
  wire  _T_1188 = _T_1184 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393289:6]
  wire  _T_1189 = ~_T_1188; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393290:6]
  wire [7:0] c_size_lookup = _c_size_lookup_T_7[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 393143:4 Monitor.scala 747:21 chipyard.TestHarness.SmallBoomConfig.fir 393162:4]
  wire  _T_1194 = _GEN_80 == c_size_lookup; // @[Monitor.scala 795:36 chipyard.TestHarness.SmallBoomConfig.fir 393308:8]
  wire  _T_1196 = _T_1194 | reset; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393310:8]
  wire  _T_1197 = ~_T_1196; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393311:8]
  wire [7:0] d_sizes_clr_1 = _GEN_69[7:0]; // @[chipyard.TestHarness.SmallBoomConfig.fir 393236:4]
  wire [7:0] _inflight_sizes_T_4 = ~d_sizes_clr_1; // @[Monitor.scala 811:58 chipyard.TestHarness.SmallBoomConfig.fir 393361:4]
  wire [7:0] _inflight_sizes_T_5 = inflight_sizes_1 & _inflight_sizes_T_4; // @[Monitor.scala 811:56 chipyard.TestHarness.SmallBoomConfig.fir 393362:4]
  wire  _GEN_90 = io_in_a_valid & _T_15; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391291:10]
  wire  _GEN_100 = io_in_a_valid & _T_171; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391481:10]
  wire  _GEN_112 = io_in_a_valid & _T_331; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391619:10]
  wire  _GEN_120 = io_in_a_valid & _T_426; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391811:10]
  wire  _GEN_126 = io_in_a_valid & _T_517; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391924:10]
  wire  _GEN_132 = io_in_a_valid & _T_610; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392034:10]
  wire  _GEN_138 = io_in_a_valid & _T_696; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392142:10]
  wire  _GEN_144 = io_in_a_valid & _T_782; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392255:10]
  wire  _GEN_150 = io_in_d_valid & _T_881; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392318:10]
  wire  _GEN_160 = io_in_d_valid & _T_901; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392360:10]
  wire  _GEN_170 = io_in_d_valid & _T_929; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392418:10]
  wire  _GEN_180 = io_in_d_valid & _T_958; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392477:10]
  wire  _GEN_186 = io_in_d_valid & _T_975; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392512:10]
  wire  _GEN_192 = io_in_d_valid & _T_993; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392548:10]
  wire  _GEN_198 = _T_1088 & same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392981:10]
  wire  _GEN_203 = _T_1088 & ~same_cycle_resp; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393003:10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393058:4]
    .out(plusarg_reader_out)
  );
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 393365:4]
    .out(plusarg_reader_1_out)
  );
  always @(posedge clock) begin
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392617:4]
      a_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392617:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392627:4]
      if (a_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392628:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392616:4]
          a_first_counter <= a_first_beats1_decode;
        end else begin
          a_first_counter <= 9'h0;
        end
      end else begin
        a_first_counter <= a_first_counter1;
      end
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 392682:4]
      opcode <= io_in_a_bits_opcode; // @[Monitor.scala 397:15 chipyard.TestHarness.SmallBoomConfig.fir 392683:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 392682:4]
      size <= io_in_a_bits_size; // @[Monitor.scala 399:15 chipyard.TestHarness.SmallBoomConfig.fir 392685:6]
    end
    if (_T_1045) begin // @[Monitor.scala 396:32 chipyard.TestHarness.SmallBoomConfig.fir 392682:4]
      address <= io_in_a_bits_address; // @[Monitor.scala 401:15 chipyard.TestHarness.SmallBoomConfig.fir 392687:6]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392697:4]
      d_first_counter <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392697:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392707:4]
      if (d_first) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392708:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392696:4]
          d_first_counter <= d_first_beats1_decode;
        end else begin
          d_first_counter <= 9'h0;
        end
      end else begin
        d_first_counter <= d_first_counter1;
      end
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392771:4]
      opcode_1 <= io_in_d_bits_opcode; // @[Monitor.scala 550:15 chipyard.TestHarness.SmallBoomConfig.fir 392772:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392771:4]
      param_1 <= io_in_d_bits_param; // @[Monitor.scala 551:15 chipyard.TestHarness.SmallBoomConfig.fir 392773:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392771:4]
      size_1 <= io_in_d_bits_size; // @[Monitor.scala 552:15 chipyard.TestHarness.SmallBoomConfig.fir 392774:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392771:4]
      source_1 <= io_in_d_bits_source; // @[Monitor.scala 553:15 chipyard.TestHarness.SmallBoomConfig.fir 392775:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392771:4]
      sink <= io_in_d_bits_sink; // @[Monitor.scala 554:15 chipyard.TestHarness.SmallBoomConfig.fir 392776:6]
    end
    if (_T_1073) begin // @[Monitor.scala 549:32 chipyard.TestHarness.SmallBoomConfig.fir 392771:4]
      denied <= io_in_d_bits_denied; // @[Monitor.scala 555:15 chipyard.TestHarness.SmallBoomConfig.fir 392777:6]
    end
    if (reset) begin // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 392779:4]
      inflight <= 1'h0; // @[Monitor.scala 611:27 chipyard.TestHarness.SmallBoomConfig.fir 392779:4]
    end else begin
      inflight <= _inflight_T_2; // @[Monitor.scala 702:14 chipyard.TestHarness.SmallBoomConfig.fir 393048:4]
    end
    if (reset) begin // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 392780:4]
      inflight_opcodes <= 4'h0; // @[Monitor.scala 613:35 chipyard.TestHarness.SmallBoomConfig.fir 392780:4]
    end else begin
      inflight_opcodes <= _inflight_opcodes_T_2; // @[Monitor.scala 703:22 chipyard.TestHarness.SmallBoomConfig.fir 393052:4]
    end
    if (reset) begin // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 392781:4]
      inflight_sizes <= 8'h0; // @[Monitor.scala 615:33 chipyard.TestHarness.SmallBoomConfig.fir 392781:4]
    end else begin
      inflight_sizes <= _inflight_sizes_T_2; // @[Monitor.scala 704:20 chipyard.TestHarness.SmallBoomConfig.fir 393056:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392791:4]
      a_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392791:4]
    end else if (_a_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392801:4]
      if (a_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392802:6]
        if (a_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392616:4]
          a_first_counter_1 <= a_first_beats1_decode;
        end else begin
          a_first_counter_1 <= 9'h0;
        end
      end else begin
        a_first_counter_1 <= a_first_counter1_1;
      end
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392813:4]
      d_first_counter_1 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 392813:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 392823:4]
      if (d_first_1) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 392824:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392696:4]
          d_first_counter_1 <= d_first_beats1_decode;
        end else begin
          d_first_counter_1 <= 9'h0;
        end
      end else begin
        d_first_counter_1 <= d_first_counter1_1;
      end
    end
    if (reset) begin // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 393057:4]
      watchdog <= 32'h0; // @[Monitor.scala 706:27 chipyard.TestHarness.SmallBoomConfig.fir 393057:4]
    end else if (_T_1156) begin // @[Monitor.scala 712:47 chipyard.TestHarness.SmallBoomConfig.fir 393079:4]
      watchdog <= 32'h0; // @[Monitor.scala 712:58 chipyard.TestHarness.SmallBoomConfig.fir 393080:6]
    end else begin
      watchdog <= _watchdog_T_1; // @[Monitor.scala 711:14 chipyard.TestHarness.SmallBoomConfig.fir 393075:4]
    end
    if (reset) begin // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 393084:4]
      inflight_sizes_1 <= 8'h0; // @[Monitor.scala 725:35 chipyard.TestHarness.SmallBoomConfig.fir 393084:4]
    end else begin
      inflight_sizes_1 <= _inflight_sizes_T_5; // @[Monitor.scala 811:22 chipyard.TestHarness.SmallBoomConfig.fir 393363:4]
    end
    if (reset) begin // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 393119:4]
      d_first_counter_2 <= 9'h0; // @[Edges.scala 228:27 chipyard.TestHarness.SmallBoomConfig.fir 393119:4]
    end else if (_d_first_T) begin // @[Edges.scala 234:17 chipyard.TestHarness.SmallBoomConfig.fir 393129:4]
      if (d_first_2) begin // @[Edges.scala 235:21 chipyard.TestHarness.SmallBoomConfig.fir 393130:6]
        if (d_first_beats1_opdata) begin // @[Edges.scala 220:14 chipyard.TestHarness.SmallBoomConfig.fir 392696:4]
          d_first_counter_2 <= d_first_beats1_decode;
        end else begin
          d_first_counter_2 <= 9'h0;
        end
      end else begin
        d_first_counter_2 <= d_first_counter1_2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_15 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391291:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391292:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391358:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391359:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391373:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391374:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391380:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391381:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391397:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_90 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391398:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_171 & _T_84) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391481:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_84) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391482:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391548:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391549:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391563:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_154) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391564:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391570:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391571:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391586:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_147) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391587:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391595:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_100 & _T_166) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391596:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_331 & _T_340) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391619:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_340) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391620:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391690:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_407) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391691:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391704:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391705:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Get contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391720:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_112 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391721:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_426 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391811:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391812:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391825:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391826:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutFull contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391841:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_120 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391842:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_517 & _T_502) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391924:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_502) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391925:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391938:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391939:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel PutPartial contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391956:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_126 & _T_609) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 391957:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_610 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392034:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392035:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392048:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392049:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392064:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_132 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392065:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_696 & _T_681) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392142:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_681) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392143:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392156:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392157:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Logical contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392172:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_138 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392173:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_a_valid & _T_782 & _T_858) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392255:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_858) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392256:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint address not aligned to size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392269:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_157) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392270:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel Hint contains invalid mask (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392285:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_144 & _T_421) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392286:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel has invalid opcode (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392304:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_880) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392305:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_881 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392318:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392319:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392326:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392327:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392334:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392335:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392342:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392343:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel ReleaseAck is denied (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392350:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_150 & _T_900) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392351:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_901 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392360:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392361:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392375:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392376:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392383:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392384:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392391:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392392:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel Grant is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392399:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_160 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392400:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_929 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392418:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392419:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData smaller than a beat (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392433:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_888) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392434:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries invalid cap param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392441:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_915) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392442:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData carries toN param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392449:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_919) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392450:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392458:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_170 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392459:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_958 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392477:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392478:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392485:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392486:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392493:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_180 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392494:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_975 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392512:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392513:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392520:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392521:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392529:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_186 & _T_952) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392530:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_993 & _T_884) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392548:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_884) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392549:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck carries invalid param (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392556:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_892) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392557:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel HintAck is corrupt (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392564:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_192 & _T_896) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392565:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392644:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1027) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392645:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392660:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1035) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392661:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel address changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392676:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1023 & _T_1043) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392677:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel opcode changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392725:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1051) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392726:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel param changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392733:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1055) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392734:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel size changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392741:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1059) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392742:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel source changed within multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392749:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1063) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392750:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel sink changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392757:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1067) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392758:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel denied changed with multibeat operation (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392765:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1047 & _T_1071) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392766:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' channel re-used a source ID (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392910:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1077 & _T_1084) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 392911:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392970:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1088 & _T_1103) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392971:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & same_cycle_resp & _T_1109) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392981:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1109) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392982:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392989:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_198 & _T_1113) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 392990:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1088 & ~same_cycle_resp & _T_1121) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper opcode response (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393003:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1121) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393004:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393011:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_203 & _T_1125) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393012:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fwrite(32'h80000002,"Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n"); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393030:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1132 & _T_1137) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393031:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1144) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'A' and 'D' concurrent, despite minlatency 8 (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393042:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1144) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393043:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1153) begin
          $fwrite(32'h80000002,
            "Assertion failed: TileLink timeout expired (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:42 assert(cond, message)\n"
            ); // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393070:6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1153) begin
          $fatal; // @[Monitor.scala 42:11 chipyard.TestHarness.SmallBoomConfig.fir 393071:6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel acknowledged for nothing inflight (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393292:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1189) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393293:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fwrite(32'h80000002,
            "Assertion failed: 'D' channel contains improper response size (connected at SerialAdapter.scala:331:39)\n    at Monitor.scala:49 assert(cond, message)\n"
            ); // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393313:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1176 & _T_1197) begin
          $fatal; // @[Monitor.scala 49:11 chipyard.TestHarness.SmallBoomConfig.fir 393314:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  a_first_counter = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  address = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  d_first_counter = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  opcode_1 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  param_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  size_1 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  source_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sink = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  denied = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inflight = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  inflight_opcodes = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  inflight_sizes = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  a_first_counter_1 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  d_first_counter_1 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  watchdog = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  inflight_sizes_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  d_first_counter_2 = _RAND_18[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLBuffer_21_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393520:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393521:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393522:4]
  output        auto_in_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input         auto_in_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [2:0]  auto_in_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [3:0]  auto_in_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [31:0] auto_in_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [7:0]  auto_in_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [63:0] auto_in_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input         auto_in_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output        auto_in_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output [63:0] auto_in_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input         auto_out_a_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output        auto_out_a_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output [2:0]  auto_out_a_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output [2:0]  auto_out_a_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output [3:0]  auto_out_a_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output        auto_out_a_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output [31:0] auto_out_a_bits_address, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output [7:0]  auto_out_a_bits_mask, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output [63:0] auto_out_a_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output        auto_out_a_bits_corrupt, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  output        auto_out_d_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input         auto_out_d_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [2:0]  auto_out_d_bits_opcode, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [1:0]  auto_out_d_bits_param, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [3:0]  auto_out_d_bits_size, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input         auto_out_d_bits_source, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [2:0]  auto_out_d_bits_sink, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input         auto_out_d_bits_denied, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input  [63:0] auto_out_d_bits_data, // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
  input         auto_out_d_bits_corrupt // @[chipyard.TestHarness.SmallBoomConfig.fir 393523:4]
);
  wire  monitor_clock; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_reset; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_io_in_a_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_io_in_a_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [2:0] monitor_io_in_a_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [3:0] monitor_io_in_a_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [31:0] monitor_io_in_a_bits_address; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [7:0] monitor_io_in_a_bits_mask; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_io_in_d_ready; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_io_in_d_valid; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [2:0] monitor_io_in_d_bits_opcode; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [1:0] monitor_io_in_d_bits_param; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [3:0] monitor_io_in_d_bits_size; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_io_in_d_bits_source; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire [2:0] monitor_io_in_d_bits_sink; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_io_in_d_bits_denied; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  monitor_io_in_d_bits_corrupt; // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
  wire  bundleOut_0_a_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleOut_0_a_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleOut_0_a_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleOut_0_a_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [2:0] bundleOut_0_a_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [3:0] bundleOut_0_a_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [31:0] bundleOut_0_a_q_io_enq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [7:0] bundleOut_0_a_q_io_enq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [63:0] bundleOut_0_a_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleOut_0_a_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleOut_0_a_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [2:0] bundleOut_0_a_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [3:0] bundleOut_0_a_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleOut_0_a_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [31:0] bundleOut_0_a_q_io_deq_bits_address; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [7:0] bundleOut_0_a_q_io_deq_bits_mask; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire [63:0] bundleOut_0_a_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleOut_0_a_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
  wire  bundleIn_0_d_q_clock; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_reset; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_enq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_enq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [1:0] bundleIn_0_d_q_io_enq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [3:0] bundleIn_0_d_q_io_enq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_enq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [2:0] bundleIn_0_d_q_io_enq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_enq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [63:0] bundleIn_0_d_q_io_enq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_enq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_deq_ready; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_deq_valid; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_opcode; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [1:0] bundleIn_0_d_q_io_deq_bits_param; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [3:0] bundleIn_0_d_q_io_deq_bits_size; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_deq_bits_source; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [2:0] bundleIn_0_d_q_io_deq_bits_sink; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_deq_bits_denied; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire [63:0] bundleIn_0_d_q_io_deq_bits_data; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  wire  bundleIn_0_d_q_io_deq_bits_corrupt; // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
  TLMonitor_57_inTestHarness monitor ( // @[Nodes.scala 24:25 chipyard.TestHarness.SmallBoomConfig.fir 393530:4]
    .clock(monitor_clock),
    .reset(monitor_reset),
    .io_in_a_ready(monitor_io_in_a_ready),
    .io_in_a_valid(monitor_io_in_a_valid),
    .io_in_a_bits_opcode(monitor_io_in_a_bits_opcode),
    .io_in_a_bits_size(monitor_io_in_a_bits_size),
    .io_in_a_bits_address(monitor_io_in_a_bits_address),
    .io_in_a_bits_mask(monitor_io_in_a_bits_mask),
    .io_in_d_ready(monitor_io_in_d_ready),
    .io_in_d_valid(monitor_io_in_d_valid),
    .io_in_d_bits_opcode(monitor_io_in_d_bits_opcode),
    .io_in_d_bits_param(monitor_io_in_d_bits_param),
    .io_in_d_bits_size(monitor_io_in_d_bits_size),
    .io_in_d_bits_source(monitor_io_in_d_bits_source),
    .io_in_d_bits_sink(monitor_io_in_d_bits_sink),
    .io_in_d_bits_denied(monitor_io_in_d_bits_denied),
    .io_in_d_bits_corrupt(monitor_io_in_d_bits_corrupt)
  );
  Queue_6_inTestHarness bundleOut_0_a_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393557:4]
    .clock(bundleOut_0_a_q_clock),
    .reset(bundleOut_0_a_q_reset),
    .io_enq_ready(bundleOut_0_a_q_io_enq_ready),
    .io_enq_valid(bundleOut_0_a_q_io_enq_valid),
    .io_enq_bits_opcode(bundleOut_0_a_q_io_enq_bits_opcode),
    .io_enq_bits_size(bundleOut_0_a_q_io_enq_bits_size),
    .io_enq_bits_address(bundleOut_0_a_q_io_enq_bits_address),
    .io_enq_bits_mask(bundleOut_0_a_q_io_enq_bits_mask),
    .io_enq_bits_data(bundleOut_0_a_q_io_enq_bits_data),
    .io_deq_ready(bundleOut_0_a_q_io_deq_ready),
    .io_deq_valid(bundleOut_0_a_q_io_deq_valid),
    .io_deq_bits_opcode(bundleOut_0_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleOut_0_a_q_io_deq_bits_param),
    .io_deq_bits_size(bundleOut_0_a_q_io_deq_bits_size),
    .io_deq_bits_source(bundleOut_0_a_q_io_deq_bits_source),
    .io_deq_bits_address(bundleOut_0_a_q_io_deq_bits_address),
    .io_deq_bits_mask(bundleOut_0_a_q_io_deq_bits_mask),
    .io_deq_bits_data(bundleOut_0_a_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleOut_0_a_q_io_deq_bits_corrupt)
  );
  Queue_7_inTestHarness bundleIn_0_d_q ( // @[Decoupled.scala 296:21 chipyard.TestHarness.SmallBoomConfig.fir 393571:4]
    .clock(bundleIn_0_d_q_clock),
    .reset(bundleIn_0_d_q_reset),
    .io_enq_ready(bundleIn_0_d_q_io_enq_ready),
    .io_enq_valid(bundleIn_0_d_q_io_enq_valid),
    .io_enq_bits_opcode(bundleIn_0_d_q_io_enq_bits_opcode),
    .io_enq_bits_param(bundleIn_0_d_q_io_enq_bits_param),
    .io_enq_bits_size(bundleIn_0_d_q_io_enq_bits_size),
    .io_enq_bits_source(bundleIn_0_d_q_io_enq_bits_source),
    .io_enq_bits_sink(bundleIn_0_d_q_io_enq_bits_sink),
    .io_enq_bits_denied(bundleIn_0_d_q_io_enq_bits_denied),
    .io_enq_bits_data(bundleIn_0_d_q_io_enq_bits_data),
    .io_enq_bits_corrupt(bundleIn_0_d_q_io_enq_bits_corrupt),
    .io_deq_ready(bundleIn_0_d_q_io_deq_ready),
    .io_deq_valid(bundleIn_0_d_q_io_deq_valid),
    .io_deq_bits_opcode(bundleIn_0_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(bundleIn_0_d_q_io_deq_bits_param),
    .io_deq_bits_size(bundleIn_0_d_q_io_deq_bits_size),
    .io_deq_bits_source(bundleIn_0_d_q_io_deq_bits_source),
    .io_deq_bits_sink(bundleIn_0_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(bundleIn_0_d_q_io_deq_bits_denied),
    .io_deq_bits_data(bundleIn_0_d_q_io_deq_bits_data),
    .io_deq_bits_corrupt(bundleIn_0_d_q_io_deq_bits_corrupt)
  );
  assign auto_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 393569:4]
  assign auto_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign auto_in_d_bits_data = bundleIn_0_d_q_io_deq_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign auto_out_a_valid = bundleOut_0_a_q_io_deq_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_opcode = bundleOut_0_a_q_io_deq_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_param = bundleOut_0_a_q_io_deq_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_size = bundleOut_0_a_q_io_deq_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_source = bundleOut_0_a_q_io_deq_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_address = bundleOut_0_a_q_io_deq_bits_address; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_mask = bundleOut_0_a_q_io_deq_bits_mask; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_data = bundleOut_0_a_q_io_deq_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_a_bits_corrupt = bundleOut_0_a_q_io_deq_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Buffer.scala 37:13 chipyard.TestHarness.SmallBoomConfig.fir 393570:4]
  assign auto_out_d_ready = bundleIn_0_d_q_io_enq_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 393583:4]
  assign monitor_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393531:4]
  assign monitor_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393532:4]
  assign monitor_io_in_a_ready = bundleOut_0_a_q_io_enq_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Decoupled.scala 299:17 chipyard.TestHarness.SmallBoomConfig.fir 393569:4]
  assign monitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign monitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign monitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign monitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign monitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign monitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign monitor_io_in_d_valid = bundleIn_0_d_q_io_deq_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign monitor_io_in_d_bits_opcode = bundleIn_0_d_q_io_deq_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign monitor_io_in_d_bits_param = bundleIn_0_d_q_io_deq_bits_param; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign monitor_io_in_d_bits_size = bundleIn_0_d_q_io_deq_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign monitor_io_in_d_bits_source = bundleIn_0_d_q_io_deq_bits_source; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign monitor_io_in_d_bits_sink = bundleIn_0_d_q_io_deq_bits_sink; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign monitor_io_in_d_bits_denied = bundleIn_0_d_q_io_deq_bits_denied; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign monitor_io_in_d_bits_corrupt = bundleIn_0_d_q_io_deq_bits_corrupt; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 Buffer.scala 38:13 chipyard.TestHarness.SmallBoomConfig.fir 393584:4]
  assign bundleOut_0_a_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393558:4]
  assign bundleOut_0_a_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393559:4]
  assign bundleOut_0_a_q_io_enq_valid = auto_in_a_valid; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign bundleOut_0_a_q_io_enq_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign bundleOut_0_a_q_io_enq_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign bundleOut_0_a_q_io_enq_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign bundleOut_0_a_q_io_enq_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign bundleOut_0_a_q_io_enq_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
  assign bundleOut_0_a_q_io_deq_ready = auto_out_a_ready; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393572:4]
  assign bundleIn_0_d_q_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393573:4]
  assign bundleIn_0_d_q_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_param = auto_out_d_bits_param; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_denied = auto_out_d_bits_denied; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_enq_bits_corrupt = auto_out_d_bits_corrupt; // @[Nodes.scala 1207:84 chipyard.TestHarness.SmallBoomConfig.fir 393553:4 LazyModule.scala 311:12 chipyard.TestHarness.SmallBoomConfig.fir 393555:4]
  assign bundleIn_0_d_q_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1210:84 chipyard.TestHarness.SmallBoomConfig.fir 393528:4 LazyModule.scala 309:16 chipyard.TestHarness.SmallBoomConfig.fir 393556:4]
endmodule




module SerialRAM_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393604:2]
  input         clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393605:4]
  input         reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393606:4]
  input         io_ser_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  output        io_ser_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  output [3:0]  io_ser_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  output        io_ser_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  input         io_ser_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  input  [3:0]  io_ser_out_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  output        io_tsi_ser_in_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  input         io_tsi_ser_in_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  input  [31:0] io_tsi_ser_in_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  input         io_tsi_ser_out_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  output        io_tsi_ser_out_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
  output [31:0] io_tsi_ser_out_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 393608:4]
);
  wire  adapter_clock; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_reset; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_auto_out_a_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_auto_out_a_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [2:0] adapter_auto_out_a_bits_opcode; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [3:0] adapter_auto_out_a_bits_size; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [31:0] adapter_auto_out_a_bits_address; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [7:0] adapter_auto_out_a_bits_mask; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [63:0] adapter_auto_out_a_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_auto_out_d_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_auto_out_d_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [63:0] adapter_auto_out_d_bits_data; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_io_serial_in_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_io_serial_in_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [31:0] adapter_io_serial_in_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_io_serial_out_ready; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  adapter_io_serial_out_valid; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire [31:0] adapter_io_serial_out_bits; // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
  wire  serdesser_clock; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_reset; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_manager_in_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [3:0] serdesser_auto_manager_in_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [31:0] serdesser_auto_manager_in_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [7:0] serdesser_auto_manager_in_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [63:0] serdesser_auto_manager_in_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [1:0] serdesser_auto_manager_in_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [3:0] serdesser_auto_manager_in_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_manager_in_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [63:0] serdesser_auto_manager_in_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_manager_in_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_a_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_a_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_client_out_a_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_client_out_a_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_client_out_a_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [3:0] serdesser_auto_client_out_a_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [28:0] serdesser_auto_client_out_a_bits_address; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [7:0] serdesser_auto_client_out_a_bits_mask; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [63:0] serdesser_auto_client_out_a_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_a_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_d_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_d_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_client_out_d_bits_opcode; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [1:0] serdesser_auto_client_out_d_bits_param; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [2:0] serdesser_auto_client_out_d_bits_size; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [3:0] serdesser_auto_client_out_d_bits_source; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_d_bits_sink; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_d_bits_denied; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [63:0] serdesser_auto_client_out_d_bits_data; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_auto_client_out_d_bits_corrupt; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_io_ser_in_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_io_ser_in_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [3:0] serdesser_io_ser_in_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_io_ser_out_ready; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  serdesser_io_ser_out_valid; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire [3:0] serdesser_io_ser_out_bits; // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
  wire  srams_clock; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire  srams_reset; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire  srams_auto_in_a_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire  srams_auto_in_a_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [2:0] srams_auto_in_a_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [2:0] srams_auto_in_a_bits_param; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [1:0] srams_auto_in_a_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [7:0] srams_auto_in_a_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [28:0] srams_auto_in_a_bits_address; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [7:0] srams_auto_in_a_bits_mask; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [63:0] srams_auto_in_a_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire  srams_auto_in_a_bits_corrupt; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire  srams_auto_in_d_ready; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire  srams_auto_in_d_valid; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [2:0] srams_auto_in_d_bits_opcode; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [1:0] srams_auto_in_d_bits_size; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [7:0] srams_auto_in_d_bits_source; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire [63:0] srams_auto_in_d_bits_data; // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
  wire  xbar_auto_in_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_in_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_in_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_in_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_in_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [3:0] xbar_auto_in_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [28:0] xbar_auto_in_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [7:0] xbar_auto_in_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [63:0] xbar_auto_in_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_in_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_in_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_in_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_in_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [1:0] xbar_auto_in_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_in_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [3:0] xbar_auto_in_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_in_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_in_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [63:0] xbar_auto_in_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_in_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_a_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_a_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_out_a_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_out_a_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [3:0] xbar_auto_out_a_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [28:0] xbar_auto_out_a_bits_address; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [7:0] xbar_auto_out_a_bits_mask; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [63:0] xbar_auto_out_a_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_a_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_d_ready; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_d_valid; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [1:0] xbar_auto_out_d_bits_param; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [2:0] xbar_auto_out_d_bits_size; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [3:0] xbar_auto_out_d_bits_source; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_d_bits_sink; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_d_bits_denied; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire [63:0] xbar_auto_out_d_bits_data; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  xbar_auto_out_d_bits_corrupt; // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
  wire  buffer_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [2:0] buffer_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [2:0] buffer_auto_in_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [1:0] buffer_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [7:0] buffer_auto_in_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [28:0] buffer_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [7:0] buffer_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [63:0] buffer_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [2:0] buffer_auto_in_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [1:0] buffer_auto_in_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [1:0] buffer_auto_in_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [7:0] buffer_auto_in_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [63:0] buffer_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_in_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [2:0] buffer_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [2:0] buffer_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [1:0] buffer_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [7:0] buffer_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [28:0] buffer_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [7:0] buffer_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [63:0] buffer_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  buffer_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [2:0] buffer_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [1:0] buffer_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [7:0] buffer_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire [63:0] buffer_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
  wire  fragmenter_clock; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_reset; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_in_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_in_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_in_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [3:0] fragmenter_auto_in_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [28:0] fragmenter_auto_in_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [7:0] fragmenter_auto_in_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [63:0] fragmenter_auto_in_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_in_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [1:0] fragmenter_auto_in_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_in_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [3:0] fragmenter_auto_in_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [63:0] fragmenter_auto_in_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_in_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_a_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_a_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_out_a_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_out_a_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [1:0] fragmenter_auto_out_a_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [7:0] fragmenter_auto_out_a_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [28:0] fragmenter_auto_out_a_bits_address; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [7:0] fragmenter_auto_out_a_bits_mask; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [63:0] fragmenter_auto_out_a_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_a_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_d_ready; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_d_valid; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [2:0] fragmenter_auto_out_d_bits_opcode; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [1:0] fragmenter_auto_out_d_bits_param; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [1:0] fragmenter_auto_out_d_bits_size; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [7:0] fragmenter_auto_out_d_bits_source; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_d_bits_sink; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_d_bits_denied; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire [63:0] fragmenter_auto_out_d_bits_data; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  fragmenter_auto_out_d_bits_corrupt; // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
  wire  buffer_1_clock; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_reset; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_in_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_in_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [2:0] buffer_1_auto_in_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [3:0] buffer_1_auto_in_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [31:0] buffer_1_auto_in_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [7:0] buffer_1_auto_in_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [63:0] buffer_1_auto_in_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_in_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_in_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [63:0] buffer_1_auto_in_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_a_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_a_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [2:0] buffer_1_auto_out_a_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [2:0] buffer_1_auto_out_a_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [3:0] buffer_1_auto_out_a_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_a_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [31:0] buffer_1_auto_out_a_bits_address; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [7:0] buffer_1_auto_out_a_bits_mask; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [63:0] buffer_1_auto_out_a_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_a_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_d_ready; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_d_valid; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [2:0] buffer_1_auto_out_d_bits_opcode; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [1:0] buffer_1_auto_out_d_bits_param; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [3:0] buffer_1_auto_out_d_bits_size; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_d_bits_source; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [2:0] buffer_1_auto_out_d_bits_sink; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_d_bits_denied; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire [63:0] buffer_1_auto_out_d_bits_data; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  wire  buffer_1_auto_out_d_bits_corrupt; // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
  SerialAdapter_inTestHarness adapter ( // @[SerialAdapter.scala 311:27 chipyard.TestHarness.SmallBoomConfig.fir 393614:4]
    .clock(adapter_clock),
    .reset(adapter_reset),
    .auto_out_a_ready(adapter_auto_out_a_ready),
    .auto_out_a_valid(adapter_auto_out_a_valid),
    .auto_out_a_bits_opcode(adapter_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(adapter_auto_out_a_bits_size),
    .auto_out_a_bits_address(adapter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(adapter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(adapter_auto_out_a_bits_data),
    .auto_out_d_ready(adapter_auto_out_d_ready),
    .auto_out_d_valid(adapter_auto_out_d_valid),
    .auto_out_d_bits_data(adapter_auto_out_d_bits_data),
    .io_serial_in_ready(adapter_io_serial_in_ready),
    .io_serial_in_valid(adapter_io_serial_in_valid),
    .io_serial_in_bits(adapter_io_serial_in_bits),
    .io_serial_out_ready(adapter_io_serial_out_ready),
    .io_serial_out_valid(adapter_io_serial_out_valid),
    .io_serial_out_bits(adapter_io_serial_out_bits)
  );
  TLSerdesser_1_inTestHarness serdesser ( // @[SerialAdapter.scala 312:29 chipyard.TestHarness.SmallBoomConfig.fir 393621:4]
    .clock(serdesser_clock),
    .reset(serdesser_reset),
    .auto_manager_in_a_ready(serdesser_auto_manager_in_a_ready),
    .auto_manager_in_a_valid(serdesser_auto_manager_in_a_valid),
    .auto_manager_in_a_bits_opcode(serdesser_auto_manager_in_a_bits_opcode),
    .auto_manager_in_a_bits_param(serdesser_auto_manager_in_a_bits_param),
    .auto_manager_in_a_bits_size(serdesser_auto_manager_in_a_bits_size),
    .auto_manager_in_a_bits_source(serdesser_auto_manager_in_a_bits_source),
    .auto_manager_in_a_bits_address(serdesser_auto_manager_in_a_bits_address),
    .auto_manager_in_a_bits_mask(serdesser_auto_manager_in_a_bits_mask),
    .auto_manager_in_a_bits_data(serdesser_auto_manager_in_a_bits_data),
    .auto_manager_in_a_bits_corrupt(serdesser_auto_manager_in_a_bits_corrupt),
    .auto_manager_in_d_ready(serdesser_auto_manager_in_d_ready),
    .auto_manager_in_d_valid(serdesser_auto_manager_in_d_valid),
    .auto_manager_in_d_bits_opcode(serdesser_auto_manager_in_d_bits_opcode),
    .auto_manager_in_d_bits_param(serdesser_auto_manager_in_d_bits_param),
    .auto_manager_in_d_bits_size(serdesser_auto_manager_in_d_bits_size),
    .auto_manager_in_d_bits_source(serdesser_auto_manager_in_d_bits_source),
    .auto_manager_in_d_bits_sink(serdesser_auto_manager_in_d_bits_sink),
    .auto_manager_in_d_bits_denied(serdesser_auto_manager_in_d_bits_denied),
    .auto_manager_in_d_bits_data(serdesser_auto_manager_in_d_bits_data),
    .auto_manager_in_d_bits_corrupt(serdesser_auto_manager_in_d_bits_corrupt),
    .auto_client_out_a_ready(serdesser_auto_client_out_a_ready),
    .auto_client_out_a_valid(serdesser_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(serdesser_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_param(serdesser_auto_client_out_a_bits_param),
    .auto_client_out_a_bits_size(serdesser_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(serdesser_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(serdesser_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(serdesser_auto_client_out_a_bits_mask),
    .auto_client_out_a_bits_data(serdesser_auto_client_out_a_bits_data),
    .auto_client_out_a_bits_corrupt(serdesser_auto_client_out_a_bits_corrupt),
    .auto_client_out_d_ready(serdesser_auto_client_out_d_ready),
    .auto_client_out_d_valid(serdesser_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(serdesser_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_param(serdesser_auto_client_out_d_bits_param),
    .auto_client_out_d_bits_size(serdesser_auto_client_out_d_bits_size),
    .auto_client_out_d_bits_source(serdesser_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_sink(serdesser_auto_client_out_d_bits_sink),
    .auto_client_out_d_bits_denied(serdesser_auto_client_out_d_bits_denied),
    .auto_client_out_d_bits_data(serdesser_auto_client_out_d_bits_data),
    .auto_client_out_d_bits_corrupt(serdesser_auto_client_out_d_bits_corrupt),
    .io_ser_in_ready(serdesser_io_ser_in_ready),
    .io_ser_in_valid(serdesser_io_ser_in_valid),
    .io_ser_in_bits(serdesser_io_ser_in_bits),
    .io_ser_out_ready(serdesser_io_ser_out_ready),
    .io_ser_out_valid(serdesser_io_ser_out_valid),
    .io_ser_out_bits(serdesser_io_ser_out_bits)
  );
  TLRAM_inTestHarness srams ( // @[SerialAdapter.scala 322:15 chipyard.TestHarness.SmallBoomConfig.fir 393628:4]
    .clock(srams_clock),
    .reset(srams_reset),
    .auto_in_a_ready(srams_auto_in_a_ready),
    .auto_in_a_valid(srams_auto_in_a_valid),
    .auto_in_a_bits_opcode(srams_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(srams_auto_in_a_bits_param),
    .auto_in_a_bits_size(srams_auto_in_a_bits_size),
    .auto_in_a_bits_source(srams_auto_in_a_bits_source),
    .auto_in_a_bits_address(srams_auto_in_a_bits_address),
    .auto_in_a_bits_mask(srams_auto_in_a_bits_mask),
    .auto_in_a_bits_data(srams_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(srams_auto_in_a_bits_corrupt),
    .auto_in_d_ready(srams_auto_in_d_ready),
    .auto_in_d_valid(srams_auto_in_d_valid),
    .auto_in_d_bits_opcode(srams_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(srams_auto_in_d_bits_size),
    .auto_in_d_bits_source(srams_auto_in_d_bits_source),
    .auto_in_d_bits_data(srams_auto_in_d_bits_data)
  );
  TLXbar_10_inTestHarness xbar ( // @[Xbar.scala 142:26 chipyard.TestHarness.SmallBoomConfig.fir 393634:4]
    .auto_in_a_ready(xbar_auto_in_a_ready),
    .auto_in_a_valid(xbar_auto_in_a_valid),
    .auto_in_a_bits_opcode(xbar_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(xbar_auto_in_a_bits_param),
    .auto_in_a_bits_size(xbar_auto_in_a_bits_size),
    .auto_in_a_bits_source(xbar_auto_in_a_bits_source),
    .auto_in_a_bits_address(xbar_auto_in_a_bits_address),
    .auto_in_a_bits_mask(xbar_auto_in_a_bits_mask),
    .auto_in_a_bits_data(xbar_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(xbar_auto_in_a_bits_corrupt),
    .auto_in_d_ready(xbar_auto_in_d_ready),
    .auto_in_d_valid(xbar_auto_in_d_valid),
    .auto_in_d_bits_opcode(xbar_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(xbar_auto_in_d_bits_param),
    .auto_in_d_bits_size(xbar_auto_in_d_bits_size),
    .auto_in_d_bits_source(xbar_auto_in_d_bits_source),
    .auto_in_d_bits_sink(xbar_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(xbar_auto_in_d_bits_denied),
    .auto_in_d_bits_data(xbar_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(xbar_auto_in_d_bits_corrupt),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(xbar_auto_out_a_bits_corrupt),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(xbar_auto_out_d_bits_param),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(xbar_auto_out_d_bits_denied),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(xbar_auto_out_d_bits_corrupt)
  );
  TLBuffer_20_inTestHarness buffer ( // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393640:4]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_a_ready(buffer_auto_in_a_ready),
    .auto_in_a_valid(buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(buffer_auto_in_a_bits_corrupt),
    .auto_in_d_ready(buffer_auto_in_d_ready),
    .auto_in_d_valid(buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(buffer_auto_in_d_bits_param),
    .auto_in_d_bits_size(buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(buffer_auto_in_d_bits_denied),
    .auto_in_d_bits_data(buffer_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(buffer_auto_in_d_bits_corrupt),
    .auto_out_a_ready(buffer_auto_out_a_ready),
    .auto_out_a_valid(buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_auto_out_d_ready),
    .auto_out_d_valid(buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_auto_out_d_bits_source),
    .auto_out_d_bits_data(buffer_auto_out_d_bits_data)
  );
  TLFragmenter_7_inTestHarness fragmenter ( // @[Fragmenter.scala 333:34 chipyard.TestHarness.SmallBoomConfig.fir 393646:4]
    .clock(fragmenter_clock),
    .reset(fragmenter_reset),
    .auto_in_a_ready(fragmenter_auto_in_a_ready),
    .auto_in_a_valid(fragmenter_auto_in_a_valid),
    .auto_in_a_bits_opcode(fragmenter_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(fragmenter_auto_in_a_bits_param),
    .auto_in_a_bits_size(fragmenter_auto_in_a_bits_size),
    .auto_in_a_bits_source(fragmenter_auto_in_a_bits_source),
    .auto_in_a_bits_address(fragmenter_auto_in_a_bits_address),
    .auto_in_a_bits_mask(fragmenter_auto_in_a_bits_mask),
    .auto_in_a_bits_data(fragmenter_auto_in_a_bits_data),
    .auto_in_a_bits_corrupt(fragmenter_auto_in_a_bits_corrupt),
    .auto_in_d_ready(fragmenter_auto_in_d_ready),
    .auto_in_d_valid(fragmenter_auto_in_d_valid),
    .auto_in_d_bits_opcode(fragmenter_auto_in_d_bits_opcode),
    .auto_in_d_bits_param(fragmenter_auto_in_d_bits_param),
    .auto_in_d_bits_size(fragmenter_auto_in_d_bits_size),
    .auto_in_d_bits_source(fragmenter_auto_in_d_bits_source),
    .auto_in_d_bits_sink(fragmenter_auto_in_d_bits_sink),
    .auto_in_d_bits_denied(fragmenter_auto_in_d_bits_denied),
    .auto_in_d_bits_data(fragmenter_auto_in_d_bits_data),
    .auto_in_d_bits_corrupt(fragmenter_auto_in_d_bits_corrupt),
    .auto_out_a_ready(fragmenter_auto_out_a_ready),
    .auto_out_a_valid(fragmenter_auto_out_a_valid),
    .auto_out_a_bits_opcode(fragmenter_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(fragmenter_auto_out_a_bits_param),
    .auto_out_a_bits_size(fragmenter_auto_out_a_bits_size),
    .auto_out_a_bits_source(fragmenter_auto_out_a_bits_source),
    .auto_out_a_bits_address(fragmenter_auto_out_a_bits_address),
    .auto_out_a_bits_mask(fragmenter_auto_out_a_bits_mask),
    .auto_out_a_bits_data(fragmenter_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(fragmenter_auto_out_a_bits_corrupt),
    .auto_out_d_ready(fragmenter_auto_out_d_ready),
    .auto_out_d_valid(fragmenter_auto_out_d_valid),
    .auto_out_d_bits_opcode(fragmenter_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(fragmenter_auto_out_d_bits_param),
    .auto_out_d_bits_size(fragmenter_auto_out_d_bits_size),
    .auto_out_d_bits_source(fragmenter_auto_out_d_bits_source),
    .auto_out_d_bits_sink(fragmenter_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(fragmenter_auto_out_d_bits_denied),
    .auto_out_d_bits_data(fragmenter_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(fragmenter_auto_out_d_bits_corrupt)
  );
  TLBuffer_21_inTestHarness buffer_1 ( // @[Buffer.scala 68:28 chipyard.TestHarness.SmallBoomConfig.fir 393652:4]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_a_ready(buffer_1_auto_in_a_ready),
    .auto_in_a_valid(buffer_1_auto_in_a_valid),
    .auto_in_a_bits_opcode(buffer_1_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(buffer_1_auto_in_a_bits_size),
    .auto_in_a_bits_address(buffer_1_auto_in_a_bits_address),
    .auto_in_a_bits_mask(buffer_1_auto_in_a_bits_mask),
    .auto_in_a_bits_data(buffer_1_auto_in_a_bits_data),
    .auto_in_d_ready(buffer_1_auto_in_d_ready),
    .auto_in_d_valid(buffer_1_auto_in_d_valid),
    .auto_in_d_bits_data(buffer_1_auto_in_d_bits_data),
    .auto_out_a_ready(buffer_1_auto_out_a_ready),
    .auto_out_a_valid(buffer_1_auto_out_a_valid),
    .auto_out_a_bits_opcode(buffer_1_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(buffer_1_auto_out_a_bits_param),
    .auto_out_a_bits_size(buffer_1_auto_out_a_bits_size),
    .auto_out_a_bits_source(buffer_1_auto_out_a_bits_source),
    .auto_out_a_bits_address(buffer_1_auto_out_a_bits_address),
    .auto_out_a_bits_mask(buffer_1_auto_out_a_bits_mask),
    .auto_out_a_bits_data(buffer_1_auto_out_a_bits_data),
    .auto_out_a_bits_corrupt(buffer_1_auto_out_a_bits_corrupt),
    .auto_out_d_ready(buffer_1_auto_out_d_ready),
    .auto_out_d_valid(buffer_1_auto_out_d_valid),
    .auto_out_d_bits_opcode(buffer_1_auto_out_d_bits_opcode),
    .auto_out_d_bits_param(buffer_1_auto_out_d_bits_param),
    .auto_out_d_bits_size(buffer_1_auto_out_d_bits_size),
    .auto_out_d_bits_source(buffer_1_auto_out_d_bits_source),
    .auto_out_d_bits_sink(buffer_1_auto_out_d_bits_sink),
    .auto_out_d_bits_denied(buffer_1_auto_out_d_bits_denied),
    .auto_out_d_bits_data(buffer_1_auto_out_d_bits_data),
    .auto_out_d_bits_corrupt(buffer_1_auto_out_d_bits_corrupt)
  );
  assign io_ser_in_valid = serdesser_io_ser_out_valid; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.SmallBoomConfig.fir 393668:4]
  assign io_ser_in_bits = serdesser_io_ser_out_bits; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.SmallBoomConfig.fir 393667:4]
  assign io_ser_out_ready = serdesser_io_ser_in_ready; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.SmallBoomConfig.fir 393666:4]
  assign io_tsi_ser_in_ready = adapter_io_serial_in_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393675:4]
  assign io_tsi_ser_out_valid = adapter_io_serial_out_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393671:4]
  assign io_tsi_ser_out_bits = adapter_io_serial_out_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393670:4]
  assign adapter_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393619:4]
  assign adapter_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393620:4]
  assign adapter_auto_out_a_ready = buffer_1_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign adapter_auto_out_d_valid = buffer_1_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign adapter_auto_out_d_bits_data = buffer_1_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign adapter_io_serial_in_valid = io_tsi_ser_in_valid; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393674:4]
  assign adapter_io_serial_in_bits = io_tsi_ser_in_bits; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393673:4]
  assign adapter_io_serial_out_ready = io_tsi_ser_out_ready; // @[SerialAdapter.scala 341:16 chipyard.TestHarness.SmallBoomConfig.fir 393672:4]
  assign serdesser_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393626:4]
  assign serdesser_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393627:4]
  assign serdesser_auto_manager_in_a_valid = buffer_1_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_opcode = buffer_1_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_param = buffer_1_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_size = buffer_1_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_source = buffer_1_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_address = buffer_1_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_mask = buffer_1_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_data = buffer_1_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_a_bits_corrupt = buffer_1_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_manager_in_d_ready = buffer_1_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign serdesser_auto_client_out_a_ready = xbar_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_valid = xbar_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_opcode = xbar_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_param = xbar_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_size = xbar_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_source = xbar_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_sink = xbar_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_denied = xbar_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_data = xbar_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_auto_client_out_d_bits_corrupt = xbar_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign serdesser_io_ser_in_valid = io_ser_out_valid; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.SmallBoomConfig.fir 393665:4]
  assign serdesser_io_ser_in_bits = io_ser_out_bits; // @[SerialAdapter.scala 339:32 chipyard.TestHarness.SmallBoomConfig.fir 393664:4]
  assign serdesser_io_ser_out_ready = io_ser_in_ready; // @[SerialAdapter.scala 340:15 chipyard.TestHarness.SmallBoomConfig.fir 393669:4]
  assign srams_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393632:4]
  assign srams_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393633:4]
  assign srams_auto_in_a_valid = buffer_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_opcode = buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_param = buffer_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_size = buffer_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_source = buffer_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_address = buffer_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_mask = buffer_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_data = buffer_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_a_bits_corrupt = buffer_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign srams_auto_in_d_ready = buffer_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign xbar_auto_in_a_valid = serdesser_auto_client_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_opcode = serdesser_auto_client_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_param = serdesser_auto_client_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_size = serdesser_auto_client_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_source = serdesser_auto_client_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_address = serdesser_auto_client_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_mask = serdesser_auto_client_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_data = serdesser_auto_client_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_a_bits_corrupt = serdesser_auto_client_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_in_d_ready = serdesser_auto_client_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393659:4]
  assign xbar_auto_out_a_ready = fragmenter_auto_in_a_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_valid = fragmenter_auto_in_d_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_opcode = fragmenter_auto_in_d_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_param = fragmenter_auto_in_d_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_size = fragmenter_auto_in_d_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_source = fragmenter_auto_in_d_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_sink = fragmenter_auto_in_d_bits_sink; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_denied = fragmenter_auto_in_d_bits_denied; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_data = fragmenter_auto_in_d_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign xbar_auto_out_d_bits_corrupt = fragmenter_auto_in_d_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign buffer_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393644:4]
  assign buffer_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393645:4]
  assign buffer_auto_in_a_valid = fragmenter_auto_out_a_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_opcode = fragmenter_auto_out_a_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_param = fragmenter_auto_out_a_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_size = fragmenter_auto_out_a_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_source = fragmenter_auto_out_a_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_address = fragmenter_auto_out_a_bits_address; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_mask = fragmenter_auto_out_a_bits_mask; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_data = fragmenter_auto_out_a_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_a_bits_corrupt = fragmenter_auto_out_a_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_in_d_ready = fragmenter_auto_out_d_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_auto_out_a_ready = srams_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign buffer_auto_out_d_valid = srams_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign buffer_auto_out_d_bits_opcode = srams_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign buffer_auto_out_d_bits_size = srams_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign buffer_auto_out_d_bits_source = srams_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign buffer_auto_out_d_bits_data = srams_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393661:4]
  assign fragmenter_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393650:4]
  assign fragmenter_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393651:4]
  assign fragmenter_auto_in_a_valid = xbar_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_param = xbar_auto_out_a_bits_param; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_size = xbar_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_source = xbar_auto_out_a_bits_source; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_address = xbar_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_mask = xbar_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_data = xbar_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_a_bits_corrupt = xbar_auto_out_a_bits_corrupt; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_in_d_ready = xbar_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393660:4]
  assign fragmenter_auto_out_a_ready = buffer_auto_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_valid = buffer_auto_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_opcode = buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_param = buffer_auto_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_size = buffer_auto_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_source = buffer_auto_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_sink = buffer_auto_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_denied = buffer_auto_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_data = buffer_auto_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign fragmenter_auto_out_d_bits_corrupt = buffer_auto_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393662:4]
  assign buffer_1_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393656:4]
  assign buffer_1_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393657:4]
  assign buffer_1_auto_in_a_valid = adapter_auto_out_a_valid; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign buffer_1_auto_in_a_bits_opcode = adapter_auto_out_a_bits_opcode; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign buffer_1_auto_in_a_bits_size = adapter_auto_out_a_bits_size; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign buffer_1_auto_in_a_bits_address = adapter_auto_out_a_bits_address; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign buffer_1_auto_in_a_bits_mask = adapter_auto_out_a_bits_mask; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign buffer_1_auto_in_a_bits_data = adapter_auto_out_a_bits_data; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign buffer_1_auto_in_d_ready = adapter_auto_out_d_ready; // @[LazyModule.scala 298:16 chipyard.TestHarness.SmallBoomConfig.fir 393658:4]
  assign buffer_1_auto_out_a_ready = serdesser_auto_manager_in_a_ready; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_valid = serdesser_auto_manager_in_d_valid; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_opcode = serdesser_auto_manager_in_d_bits_opcode; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_param = serdesser_auto_manager_in_d_bits_param; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_size = serdesser_auto_manager_in_d_bits_size; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_source = serdesser_auto_manager_in_d_bits_source; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_sink = serdesser_auto_manager_in_d_bits_sink; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_denied = serdesser_auto_manager_in_d_bits_denied; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_data = serdesser_auto_manager_in_d_bits_data; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
  assign buffer_1_auto_out_d_bits_corrupt = serdesser_auto_manager_in_d_bits_corrupt; // @[LazyModule.scala 296:16 chipyard.TestHarness.SmallBoomConfig.fir 393663:4]
endmodule
module Queue_48_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393698:2]
  input        clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393699:4]
  input        reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393700:4]
  output       io_enq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  input        io_enq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  input  [7:0] io_enq_bits, // @[chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  input        io_deq_ready, // @[chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  output       io_deq_valid, // @[chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
  output [7:0] io_deq_bits // @[chipyard.TestHarness.SmallBoomConfig.fir 393701:4]
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:127]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  wire [6:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  wire [6:0] ram_MPORT_addr; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  reg [6:0] enq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393704:4]
  reg [6:0] deq_ptr_value; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393705:4]
  reg  maybe_full; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 393706:4]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33 chipyard.TestHarness.SmallBoomConfig.fir 393707:4]
  wire  _empty_T = ~maybe_full; // @[Decoupled.scala 224:28 chipyard.TestHarness.SmallBoomConfig.fir 393708:4]
  wire  empty = ptr_match & _empty_T; // @[Decoupled.scala 224:25 chipyard.TestHarness.SmallBoomConfig.fir 393709:4]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24 chipyard.TestHarness.SmallBoomConfig.fir 393710:4]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 393711:4]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37 chipyard.TestHarness.SmallBoomConfig.fir 393714:4]
  wire [6:0] _value_T_1 = enq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393722:6]
  wire [6:0] _value_T_3 = deq_ptr_value + 7'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393728:6]
  wire  _T = do_enq != do_deq; // @[Decoupled.scala 236:16 chipyard.TestHarness.SmallBoomConfig.fir 393731:4]
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19 chipyard.TestHarness.SmallBoomConfig.fir 393737:4]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19 chipyard.TestHarness.SmallBoomConfig.fir 393735:4]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15 chipyard.TestHarness.SmallBoomConfig.fir 393740:4]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16 chipyard.TestHarness.SmallBoomConfig.fir 393703:4]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393704:4]
      enq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393704:4]
    end else if (do_enq) begin // @[Decoupled.scala 229:17 chipyard.TestHarness.SmallBoomConfig.fir 393717:4]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393723:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393705:4]
      deq_ptr_value <= 7'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393705:4]
    end else if (do_deq) begin // @[Decoupled.scala 233:17 chipyard.TestHarness.SmallBoomConfig.fir 393725:4]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393729:6]
    end
    if (reset) begin // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 393706:4]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27 chipyard.TestHarness.SmallBoomConfig.fir 393706:4]
    end else if (_T) begin // @[Decoupled.scala 236:28 chipyard.TestHarness.SmallBoomConfig.fir 393732:4]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16 chipyard.TestHarness.SmallBoomConfig.fir 393733:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UARTAdapter_inTestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393806:2]
  input   clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393807:4]
  input   reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393808:4]
  input   io_uart_txd, // @[chipyard.TestHarness.SmallBoomConfig.fir 393809:4]
  output  io_uart_rxd // @[chipyard.TestHarness.SmallBoomConfig.fir 393809:4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  txfifo_clock; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire  txfifo_reset; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire  txfifo_io_enq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire  txfifo_io_enq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire [7:0] txfifo_io_enq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire  txfifo_io_deq_ready; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire  txfifo_io_deq_valid; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire [7:0] txfifo_io_deq_bits; // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
  wire  rxfifo_clock; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire  rxfifo_reset; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire  rxfifo_io_enq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire  rxfifo_io_enq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire [7:0] rxfifo_io_enq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire  rxfifo_io_deq_ready; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire  rxfifo_io_deq_valid; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire [7:0] rxfifo_io_deq_bits; // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
  wire  sim_clock; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  wire  sim_reset; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  wire  sim_serial_in_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  wire  sim_serial_in_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  wire [7:0] sim_serial_in_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  wire  sim_serial_out_ready; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  wire  sim_serial_out_valid; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  wire [7:0] sim_serial_out_bits; // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
  reg [1:0] txState; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393817:4]
  reg [7:0] txData; // @[UARTAdapter.scala 39:19 chipyard.TestHarness.SmallBoomConfig.fir 393818:4]
  wire  _T = txState == 2'h2; // @[UARTAdapter.scala 41:49 chipyard.TestHarness.SmallBoomConfig.fir 393819:4]
  wire  _T_1 = _T & txfifo_io_enq_ready; // @[UARTAdapter.scala 41:61 chipyard.TestHarness.SmallBoomConfig.fir 393820:4]
  reg [2:0] txDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393821:4]
  wire  wrap_wrap = txDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393825:6]
  wire [2:0] _wrap_value_T_1 = txDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393827:6]
  wire  txDataWrap = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393824:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393829:6 chipyard.TestHarness.SmallBoomConfig.fir 393823:4]
  wire  _T_2 = txState == 2'h1; // @[UARTAdapter.scala 43:51 chipyard.TestHarness.SmallBoomConfig.fir 393831:4]
  wire  _T_3 = _T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 43:63 chipyard.TestHarness.SmallBoomConfig.fir 393832:4]
  reg [9:0] txBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393833:4]
  wire  wrap_wrap_1 = txBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393837:6]
  wire [9:0] _wrap_value_T_3 = txBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393839:6]
  wire  txBaudWrap = _T_3 & wrap_wrap_1; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393836:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393844:6 chipyard.TestHarness.SmallBoomConfig.fir 393835:4]
  wire  _T_4 = txState == 2'h0; // @[UARTAdapter.scala 44:53 chipyard.TestHarness.SmallBoomConfig.fir 393846:4]
  wire  _T_5 = ~io_uart_txd; // @[UARTAdapter.scala 44:80 chipyard.TestHarness.SmallBoomConfig.fir 393847:4]
  wire  _T_6 = _T_4 & _T_5; // @[UARTAdapter.scala 44:65 chipyard.TestHarness.SmallBoomConfig.fir 393848:4]
  wire  _T_7 = _T_6 & txfifo_io_enq_ready; // @[UARTAdapter.scala 44:88 chipyard.TestHarness.SmallBoomConfig.fir 393849:4]
  reg [1:0] txSlackCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393850:4]
  wire  wrap_wrap_2 = txSlackCount == 2'h3; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393854:6]
  wire [1:0] _wrap_value_T_5 = txSlackCount + 2'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393856:6]
  wire  txSlackWrap = _T_7 & wrap_wrap_2; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393853:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393858:6 chipyard.TestHarness.SmallBoomConfig.fir 393852:4]
  wire  _T_8 = 2'h0 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393860:4]
  wire  _T_9 = 2'h1 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393868:6]
  wire  _T_10 = 2'h2 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393875:8]
  wire [7:0] _GEN_35 = {{7'd0}, io_uart_txd}; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.SmallBoomConfig.fir 393878:12]
  wire [7:0] _txData_T = _GEN_35 << txDataIdx; // @[UARTAdapter.scala 60:41 chipyard.TestHarness.SmallBoomConfig.fir 393878:12]
  wire [7:0] _txData_T_1 = txData | _txData_T; // @[UARTAdapter.scala 60:26 chipyard.TestHarness.SmallBoomConfig.fir 393879:12]
  wire [1:0] _txState_T_1 = io_uart_txd ? 2'h0 : 2'h3; // @[UARTAdapter.scala 63:23 chipyard.TestHarness.SmallBoomConfig.fir 393884:12]
  wire [1:0] _GEN_11 = txfifo_io_enq_ready ? 2'h1 : txState; // @[UARTAdapter.scala 64:39 chipyard.TestHarness.SmallBoomConfig.fir 393888:12 UARTAdapter.scala 65:17 chipyard.TestHarness.SmallBoomConfig.fir 393889:14 UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393817:4]
  wire [1:0] _GEN_12 = txDataWrap ? _txState_T_1 : _GEN_11; // @[UARTAdapter.scala 62:24 chipyard.TestHarness.SmallBoomConfig.fir 393882:10 UARTAdapter.scala 63:17 chipyard.TestHarness.SmallBoomConfig.fir 393885:12]
  wire  _T_11 = 2'h3 == txState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393893:10]
  wire  _T_13 = io_uart_txd & txfifo_io_enq_ready; // @[UARTAdapter.scala 69:32 chipyard.TestHarness.SmallBoomConfig.fir 393896:12]
  wire [1:0] _GEN_13 = _T_13 ? 2'h0 : txState; // @[UARTAdapter.scala 69:56 chipyard.TestHarness.SmallBoomConfig.fir 393897:12 UARTAdapter.scala 70:17 chipyard.TestHarness.SmallBoomConfig.fir 393898:14 UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393817:4]
  wire [1:0] _GEN_14 = _T_11 ? _GEN_13 : txState; // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393894:10 UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393817:4]
  reg [1:0] rxState; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393903:4]
  reg [9:0] rxBaudCount; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393904:4]
  wire  wrap_wrap_3 = rxBaudCount == 10'h363; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393908:6]
  wire [9:0] _wrap_value_T_7 = rxBaudCount + 10'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393910:6]
  wire  rxBaudWrap = txfifo_io_enq_ready & wrap_wrap_3; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393907:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393915:6 chipyard.TestHarness.SmallBoomConfig.fir 393906:4]
  wire  _T_14 = rxState == 2'h2; // @[UARTAdapter.scala 83:49 chipyard.TestHarness.SmallBoomConfig.fir 393917:4]
  wire  _T_15 = _T_14 & txfifo_io_enq_ready; // @[UARTAdapter.scala 83:61 chipyard.TestHarness.SmallBoomConfig.fir 393918:4]
  wire  _T_16 = _T_15 & rxBaudWrap; // @[UARTAdapter.scala 83:84 chipyard.TestHarness.SmallBoomConfig.fir 393919:4]
  reg [2:0] rxDataIdx; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393920:4]
  wire  wrap_wrap_4 = rxDataIdx == 3'h7; // @[Counter.scala 72:24 chipyard.TestHarness.SmallBoomConfig.fir 393924:6]
  wire [2:0] _wrap_value_T_9 = rxDataIdx + 3'h1; // @[Counter.scala 76:24 chipyard.TestHarness.SmallBoomConfig.fir 393926:6]
  wire  rxDataWrap = _T_16 & wrap_wrap_4; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393923:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393928:6 chipyard.TestHarness.SmallBoomConfig.fir 393922:4]
  wire  _T_17 = 2'h0 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393931:4]
  wire  _T_18 = rxBaudWrap & rxfifo_io_deq_valid; // @[UARTAdapter.scala 89:24 chipyard.TestHarness.SmallBoomConfig.fir 393934:6]
  wire  _T_19 = 2'h1 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393940:6]
  wire  _T_20 = 2'h2 == rxState; // @[Conditional.scala 37:30 chipyard.TestHarness.SmallBoomConfig.fir 393948:8]
  wire [7:0] _io_uart_rxd_T = rxfifo_io_deq_bits >> rxDataIdx; // @[UARTAdapter.scala 100:42 chipyard.TestHarness.SmallBoomConfig.fir 393950:10]
  wire  _T_21 = rxDataWrap & rxBaudWrap; // @[UARTAdapter.scala 101:23 chipyard.TestHarness.SmallBoomConfig.fir 393953:10]
  wire [1:0] _GEN_28 = _T_21 ? 2'h0 : rxState; // @[UARTAdapter.scala 101:38 chipyard.TestHarness.SmallBoomConfig.fir 393954:10 UARTAdapter.scala 102:17 chipyard.TestHarness.SmallBoomConfig.fir 393955:12 UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393903:4]
  wire  _GEN_29 = _T_20 ? _io_uart_rxd_T[0] : 1'h1; // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393949:8 UARTAdapter.scala 100:19 chipyard.TestHarness.SmallBoomConfig.fir 393952:10 UARTAdapter.scala 85:15 chipyard.TestHarness.SmallBoomConfig.fir 393930:4]
  wire  _GEN_31 = _T_19 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393941:6 UARTAdapter.scala 94:19 chipyard.TestHarness.SmallBoomConfig.fir 393942:8]
  wire  _rxfifo_io_deq_ready_T_1 = _T_14 & rxDataWrap; // @[UARTAdapter.scala 106:48 chipyard.TestHarness.SmallBoomConfig.fir 393959:4]
  wire  _rxfifo_io_deq_ready_T_2 = _rxfifo_io_deq_ready_T_1 & rxBaudWrap; // @[UARTAdapter.scala 106:62 chipyard.TestHarness.SmallBoomConfig.fir 393960:4]
  Queue_48_inTestHarness txfifo ( // @[UARTAdapter.scala 32:22 chipyard.TestHarness.SmallBoomConfig.fir 393811:4]
    .clock(txfifo_clock),
    .reset(txfifo_reset),
    .io_enq_ready(txfifo_io_enq_ready),
    .io_enq_valid(txfifo_io_enq_valid),
    .io_enq_bits(txfifo_io_enq_bits),
    .io_deq_ready(txfifo_io_deq_ready),
    .io_deq_valid(txfifo_io_deq_valid),
    .io_deq_bits(txfifo_io_deq_bits)
  );
  Queue_48_inTestHarness rxfifo ( // @[UARTAdapter.scala 33:22 chipyard.TestHarness.SmallBoomConfig.fir 393814:4]
    .clock(rxfifo_clock),
    .reset(rxfifo_reset),
    .io_enq_ready(rxfifo_io_enq_ready),
    .io_enq_valid(rxfifo_io_enq_valid),
    .io_enq_bits(rxfifo_io_enq_bits),
    .io_deq_ready(rxfifo_io_deq_ready),
    .io_deq_valid(rxfifo_io_deq_valid),
    .io_deq_bits(rxfifo_io_deq_bits)
  );
  SimUART #(.UARTNO(0)) sim ( // @[UARTAdapter.scala 108:19 chipyard.TestHarness.SmallBoomConfig.fir 393963:4]
    .clock(sim_clock),
    .reset(sim_reset),
    .serial_in_ready(sim_serial_in_ready),
    .serial_in_valid(sim_serial_in_valid),
    .serial_in_bits(sim_serial_in_bits),
    .serial_out_ready(sim_serial_out_ready),
    .serial_out_valid(sim_serial_out_valid),
    .serial_out_bits(sim_serial_out_bits)
  );
  assign io_uart_rxd = _T_17 | _GEN_31; // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393932:4 UARTAdapter.scala 88:19 chipyard.TestHarness.SmallBoomConfig.fir 393933:6]
  assign txfifo_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393812:4]
  assign txfifo_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393813:4]
  assign txfifo_io_enq_valid = _T_1 & wrap_wrap; // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393824:4 Counter.scala 118:24 chipyard.TestHarness.SmallBoomConfig.fir 393829:6 chipyard.TestHarness.SmallBoomConfig.fir 393823:4]
  assign txfifo_io_enq_bits = txData; // @[UARTAdapter.scala 75:23 chipyard.TestHarness.SmallBoomConfig.fir 393901:4]
  assign txfifo_io_deq_ready = sim_serial_out_ready; // @[UARTAdapter.scala 115:23 chipyard.TestHarness.SmallBoomConfig.fir 393972:4]
  assign rxfifo_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 393815:4]
  assign rxfifo_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393816:4]
  assign rxfifo_io_enq_valid = sim_serial_in_valid; // @[UARTAdapter.scala 118:23 chipyard.TestHarness.SmallBoomConfig.fir 393974:4]
  assign rxfifo_io_enq_bits = sim_serial_in_bits; // @[UARTAdapter.scala 117:22 chipyard.TestHarness.SmallBoomConfig.fir 393973:4]
  assign rxfifo_io_deq_ready = _rxfifo_io_deq_ready_T_2 & txfifo_io_enq_ready; // @[UARTAdapter.scala 106:76 chipyard.TestHarness.SmallBoomConfig.fir 393961:4]
  assign sim_clock = clock; // @[UARTAdapter.scala 110:16 chipyard.TestHarness.SmallBoomConfig.fir 393967:4]
  assign sim_reset = reset; // @[UARTAdapter.scala 111:25 chipyard.TestHarness.SmallBoomConfig.fir 393968:4]
  assign sim_serial_in_ready = rxfifo_io_enq_ready; // @[UARTAdapter.scala 119:26 chipyard.TestHarness.SmallBoomConfig.fir 393975:4]
  assign sim_serial_out_valid = txfifo_io_deq_valid; // @[UARTAdapter.scala 114:27 chipyard.TestHarness.SmallBoomConfig.fir 393971:4]
  assign sim_serial_out_bits = txfifo_io_deq_bits; // @[UARTAdapter.scala 113:26 chipyard.TestHarness.SmallBoomConfig.fir 393970:4]
  always @(posedge clock) begin
    if (reset) begin // @[UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393817:4]
      txState <= 2'h0; // @[UARTAdapter.scala 38:24 chipyard.TestHarness.SmallBoomConfig.fir 393817:4]
    end else if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393861:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.SmallBoomConfig.fir 393862:6]
        txState <= 2'h1; // @[UARTAdapter.scala 50:17 chipyard.TestHarness.SmallBoomConfig.fir 393864:8]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393869:6]
      if (txBaudWrap) begin // @[UARTAdapter.scala 54:24 chipyard.TestHarness.SmallBoomConfig.fir 393870:8]
        txState <= 2'h2; // @[UARTAdapter.scala 55:17 chipyard.TestHarness.SmallBoomConfig.fir 393871:10]
      end
    end else if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393876:8]
      txState <= _GEN_12;
    end else begin
      txState <= _GEN_14;
    end
    if (_T_8) begin // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393861:4]
      if (txSlackWrap) begin // @[UARTAdapter.scala 48:25 chipyard.TestHarness.SmallBoomConfig.fir 393862:6]
        txData <= 8'h0; // @[UARTAdapter.scala 49:17 chipyard.TestHarness.SmallBoomConfig.fir 393863:8]
      end
    end else if (!(_T_9)) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393869:6]
      if (_T_10) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393876:8]
        if (txfifo_io_enq_ready) begin // @[UARTAdapter.scala 59:34 chipyard.TestHarness.SmallBoomConfig.fir 393877:10]
          txData <= _txData_T_1; // @[UARTAdapter.scala 60:16 chipyard.TestHarness.SmallBoomConfig.fir 393880:12]
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393821:4]
      txDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393821:4]
    end else if (_T_1) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393824:4]
      txDataIdx <= _wrap_value_T_1; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393828:6]
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393833:4]
      txBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393833:4]
    end else if (_T_3) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393836:4]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 393841:6]
        txBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 393842:8]
      end else begin
        txBaudCount <= _wrap_value_T_3; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393840:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393850:4]
      txSlackCount <= 2'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393850:4]
    end else if (_T_7) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393853:4]
      txSlackCount <= _wrap_value_T_5; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393857:6]
    end
    if (reset) begin // @[UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393903:4]
      rxState <= 2'h0; // @[UARTAdapter.scala 79:24 chipyard.TestHarness.SmallBoomConfig.fir 393903:4]
    end else if (_T_17) begin // @[Conditional.scala 40:58 chipyard.TestHarness.SmallBoomConfig.fir 393932:4]
      if (_T_18) begin // @[UARTAdapter.scala 89:48 chipyard.TestHarness.SmallBoomConfig.fir 393935:6]
        rxState <= 2'h1; // @[UARTAdapter.scala 90:17 chipyard.TestHarness.SmallBoomConfig.fir 393936:8]
      end
    end else if (_T_19) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393941:6]
      if (rxBaudWrap) begin // @[UARTAdapter.scala 95:24 chipyard.TestHarness.SmallBoomConfig.fir 393943:8]
        rxState <= 2'h2; // @[UARTAdapter.scala 96:17 chipyard.TestHarness.SmallBoomConfig.fir 393944:10]
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67 chipyard.TestHarness.SmallBoomConfig.fir 393949:8]
      rxState <= _GEN_28;
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393904:4]
      rxBaudCount <= 10'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393904:4]
    end else if (txfifo_io_enq_ready) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393907:4]
      if (wrap_wrap_3) begin // @[Counter.scala 86:20 chipyard.TestHarness.SmallBoomConfig.fir 393912:6]
        rxBaudCount <= 10'h0; // @[Counter.scala 86:28 chipyard.TestHarness.SmallBoomConfig.fir 393913:8]
      end else begin
        rxBaudCount <= _wrap_value_T_7; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393911:6]
      end
    end
    if (reset) begin // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393920:4]
      rxDataIdx <= 3'h0; // @[Counter.scala 60:40 chipyard.TestHarness.SmallBoomConfig.fir 393920:4]
    end else if (_T_16) begin // @[Counter.scala 118:17 chipyard.TestHarness.SmallBoomConfig.fir 393923:4]
      rxDataIdx <= _wrap_value_T_9; // @[Counter.scala 76:15 chipyard.TestHarness.SmallBoomConfig.fir 393927:6]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  txState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  txData = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  txDataIdx = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  txBaudCount = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  txSlackCount = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  rxState = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  rxBaudCount = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  rxDataIdx = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule


module TestHarness( // @[chipyard.TestHarness.SmallBoomConfig.fir 393977:2]
  input   clock, // @[chipyard.TestHarness.SmallBoomConfig.fir 393978:4]
  input   reset, // @[chipyard.TestHarness.SmallBoomConfig.fir 393979:4]
  output  io_success // @[chipyard.TestHarness.SmallBoomConfig.fir 393980:4]
);
  wire  chiptop_jtag_TCK; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_jtag_TMS; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_jtag_TDI; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_jtag_TDO_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_jtag_TDO_driven; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_serial_tl_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_serial_tl_bits_in_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_serial_tl_bits_in_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_serial_tl_bits_in_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_serial_tl_bits_out_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_serial_tl_bits_out_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_serial_tl_bits_out_bits; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_aw_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_aw_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [31:0] chiptop_axi4_mem_0_bits_aw_bits_addr; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [7:0] chiptop_axi4_mem_0_bits_aw_bits_len; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [2:0] chiptop_axi4_mem_0_bits_aw_bits_size; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [1:0] chiptop_axi4_mem_0_bits_aw_bits_burst; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_aw_bits_lock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_cache; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [2:0] chiptop_axi4_mem_0_bits_aw_bits_prot; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_aw_bits_qos; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_w_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_w_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [63:0] chiptop_axi4_mem_0_bits_w_bits_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [7:0] chiptop_axi4_mem_0_bits_w_bits_strb; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_w_bits_last; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_b_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_b_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_b_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [1:0] chiptop_axi4_mem_0_bits_b_bits_resp; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_ar_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_ar_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [31:0] chiptop_axi4_mem_0_bits_ar_bits_addr; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [7:0] chiptop_axi4_mem_0_bits_ar_bits_len; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [2:0] chiptop_axi4_mem_0_bits_ar_bits_size; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [1:0] chiptop_axi4_mem_0_bits_ar_bits_burst; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_ar_bits_lock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_cache; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [2:0] chiptop_axi4_mem_0_bits_ar_bits_prot; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_ar_bits_qos; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_r_ready; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_r_valid; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [3:0] chiptop_axi4_mem_0_bits_r_bits_id; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [63:0] chiptop_axi4_mem_0_bits_r_bits_data; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire [1:0] chiptop_axi4_mem_0_bits_r_bits_resp; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_axi4_mem_0_bits_r_bits_last; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_uart_0_txd; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_uart_0_rxd; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_reset_wire_reset; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  chiptop_clock; // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
  wire  SimJTAG_clock; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_reset; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_jtag_TRSTn; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_jtag_TCK; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_jtag_TMS; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_jtag_TDI; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_jtag_TDO_data; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_jtag_TDO_driven; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_enable; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire  SimJTAG_init_done; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire [31:0] SimJTAG_exit; // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 394011:4]
  wire  ram_clock; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_reset; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire [3:0] ram_io_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire [3:0] ram_io_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_tsi_ser_in_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire [31:0] ram_io_tsi_ser_in_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_tsi_ser_out_ready; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire [31:0] ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
  wire  success_sim_clock; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire  success_sim_reset; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire  success_sim_serial_in_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire  success_sim_serial_in_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire [31:0] success_sim_serial_in_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire  success_sim_serial_out_ready; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire  success_sim_serial_out_valid; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire [31:0] success_sim_serial_out_bits; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire  success_sim_exit; // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
  wire  simdram_clock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_reset; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_aw_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_aw_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_aw_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [31:0] simdram_axi_aw_bits_addr; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [7:0] simdram_axi_aw_bits_len; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [2:0] simdram_axi_aw_bits_size; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [1:0] simdram_axi_aw_bits_burst; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_aw_bits_lock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_aw_bits_cache; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [2:0] simdram_axi_aw_bits_prot; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_aw_bits_qos; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_w_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_w_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [63:0] simdram_axi_w_bits_data; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [7:0] simdram_axi_w_bits_strb; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_w_bits_last; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_b_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_b_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_b_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [1:0] simdram_axi_b_bits_resp; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_ar_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_ar_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_ar_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [31:0] simdram_axi_ar_bits_addr; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [7:0] simdram_axi_ar_bits_len; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [2:0] simdram_axi_ar_bits_size; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [1:0] simdram_axi_ar_bits_burst; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_ar_bits_lock; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_ar_bits_cache; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [2:0] simdram_axi_ar_bits_prot; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_ar_bits_qos; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_r_ready; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_r_valid; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [3:0] simdram_axi_r_bits_id; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [63:0] simdram_axi_r_bits_data; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire [1:0] simdram_axi_r_bits_resp; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  simdram_axi_r_bits_last; // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
  wire  uart_sim_0_clock; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394064:4]
  wire  uart_sim_0_reset; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394064:4]
  wire  uart_sim_0_io_uart_txd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394064:4]
  wire  uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394064:4]
  wire  dtm_success = SimJTAG_exit == 32'h1; // @[Periphery.scala 233:26 chipyard.TestHarness.SmallBoomConfig.fir 394015:4]
  wire  _T_2 = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.SmallBoomConfig.fir 394003:4]
  wire  _T_3 = SimJTAG_exit >= 32'h2; // @[Periphery.scala 234:19 chipyard.TestHarness.SmallBoomConfig.fir 394017:4]
  wire [31:0] _T_4 = {{1'd0}, SimJTAG_exit[31:1]}; // @[Periphery.scala 235:59 chipyard.TestHarness.SmallBoomConfig.fir 394019:6]

  ChipTop chiptop ( // @[TestHarness.scala 34:19 chipyard.TestHarness.SmallBoomConfig.fir 393982:4]
    .jtag_TCK(chiptop_jtag_TCK),
    .jtag_TMS(chiptop_jtag_TMS),
    .jtag_TDI(chiptop_jtag_TDI),
    .jtag_TDO_data(chiptop_jtag_TDO_data),
    .jtag_TDO_driven(chiptop_jtag_TDO_driven),
    .serial_tl_clock(chiptop_serial_tl_clock),
    .serial_tl_bits_in_ready(chiptop_serial_tl_bits_in_ready),
    .serial_tl_bits_in_valid(chiptop_serial_tl_bits_in_valid),
    .serial_tl_bits_in_bits(chiptop_serial_tl_bits_in_bits),
    .serial_tl_bits_out_ready(chiptop_serial_tl_bits_out_ready),
    .serial_tl_bits_out_valid(chiptop_serial_tl_bits_out_valid),
    .serial_tl_bits_out_bits(chiptop_serial_tl_bits_out_bits),
    .axi4_mem_0_clock(chiptop_axi4_mem_0_clock),
    .axi4_mem_0_reset(chiptop_axi4_mem_0_reset),
    .axi4_mem_0_bits_aw_ready(chiptop_axi4_mem_0_bits_aw_ready),
    .axi4_mem_0_bits_aw_valid(chiptop_axi4_mem_0_bits_aw_valid),
    .axi4_mem_0_bits_aw_bits_id(chiptop_axi4_mem_0_bits_aw_bits_id),
    .axi4_mem_0_bits_aw_bits_addr(chiptop_axi4_mem_0_bits_aw_bits_addr),
    .axi4_mem_0_bits_aw_bits_len(chiptop_axi4_mem_0_bits_aw_bits_len),
    .axi4_mem_0_bits_aw_bits_size(chiptop_axi4_mem_0_bits_aw_bits_size),
    .axi4_mem_0_bits_aw_bits_burst(chiptop_axi4_mem_0_bits_aw_bits_burst),
    .axi4_mem_0_bits_aw_bits_lock(chiptop_axi4_mem_0_bits_aw_bits_lock),
    .axi4_mem_0_bits_aw_bits_cache(chiptop_axi4_mem_0_bits_aw_bits_cache),
    .axi4_mem_0_bits_aw_bits_prot(chiptop_axi4_mem_0_bits_aw_bits_prot),
    .axi4_mem_0_bits_aw_bits_qos(chiptop_axi4_mem_0_bits_aw_bits_qos),
    .axi4_mem_0_bits_w_ready(chiptop_axi4_mem_0_bits_w_ready),
    .axi4_mem_0_bits_w_valid(chiptop_axi4_mem_0_bits_w_valid),
    .axi4_mem_0_bits_w_bits_data(chiptop_axi4_mem_0_bits_w_bits_data),
    .axi4_mem_0_bits_w_bits_strb(chiptop_axi4_mem_0_bits_w_bits_strb),
    .axi4_mem_0_bits_w_bits_last(chiptop_axi4_mem_0_bits_w_bits_last),
    .axi4_mem_0_bits_b_ready(chiptop_axi4_mem_0_bits_b_ready),
    .axi4_mem_0_bits_b_valid(chiptop_axi4_mem_0_bits_b_valid),
    .axi4_mem_0_bits_b_bits_id(chiptop_axi4_mem_0_bits_b_bits_id),
    .axi4_mem_0_bits_b_bits_resp(chiptop_axi4_mem_0_bits_b_bits_resp),
    .axi4_mem_0_bits_ar_ready(chiptop_axi4_mem_0_bits_ar_ready),
    .axi4_mem_0_bits_ar_valid(chiptop_axi4_mem_0_bits_ar_valid),
    .axi4_mem_0_bits_ar_bits_id(chiptop_axi4_mem_0_bits_ar_bits_id),
    .axi4_mem_0_bits_ar_bits_addr(chiptop_axi4_mem_0_bits_ar_bits_addr),
    .axi4_mem_0_bits_ar_bits_len(chiptop_axi4_mem_0_bits_ar_bits_len),
    .axi4_mem_0_bits_ar_bits_size(chiptop_axi4_mem_0_bits_ar_bits_size),
    .axi4_mem_0_bits_ar_bits_burst(chiptop_axi4_mem_0_bits_ar_bits_burst),
    .axi4_mem_0_bits_ar_bits_lock(chiptop_axi4_mem_0_bits_ar_bits_lock),
    .axi4_mem_0_bits_ar_bits_cache(chiptop_axi4_mem_0_bits_ar_bits_cache),
    .axi4_mem_0_bits_ar_bits_prot(chiptop_axi4_mem_0_bits_ar_bits_prot),
    .axi4_mem_0_bits_ar_bits_qos(chiptop_axi4_mem_0_bits_ar_bits_qos),
    .axi4_mem_0_bits_r_ready(chiptop_axi4_mem_0_bits_r_ready),
    .axi4_mem_0_bits_r_valid(chiptop_axi4_mem_0_bits_r_valid),
    .axi4_mem_0_bits_r_bits_id(chiptop_axi4_mem_0_bits_r_bits_id),
    .axi4_mem_0_bits_r_bits_data(chiptop_axi4_mem_0_bits_r_bits_data),
    .axi4_mem_0_bits_r_bits_resp(chiptop_axi4_mem_0_bits_r_bits_resp),
    .axi4_mem_0_bits_r_bits_last(chiptop_axi4_mem_0_bits_r_bits_last),
    .uart_0_txd(chiptop_uart_0_txd),
    .uart_0_rxd(chiptop_uart_0_rxd),
    .reset_wire_reset(chiptop_reset_wire_reset),
    .clock(chiptop_clock)
  );


  SimJTAG #(.TICK_DELAY(3)) SimJTAG ( // @[HarnessBinders.scala 190:26 chipyard.TestHarness.SmallBoomConfig.fir 393994:4]
    .clock(SimJTAG_clock),
    .reset(SimJTAG_reset),
    .jtag_TRSTn(SimJTAG_jtag_TRSTn),
    .jtag_TCK(SimJTAG_jtag_TCK),
    .jtag_TMS(SimJTAG_jtag_TMS),
    .jtag_TDI(SimJTAG_jtag_TDI),
    .jtag_TDO_data(SimJTAG_jtag_TDO_data),
    .jtag_TDO_driven(SimJTAG_jtag_TDO_driven),
    .enable(SimJTAG_enable),
    .init_done(SimJTAG_init_done),
    .exit(SimJTAG_exit)
  );


  plusarg_reader #(.FORMAT("jtag_rbb_enable=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 80:11 chipyard.TestHarness.SmallBoomConfig.fir 394011:4]
    .out(plusarg_reader_out)
  );


  SerialRAM_inTestHarness ram ( // @[SerialAdapter.scala 27:26 chipyard.TestHarness.SmallBoomConfig.fir 394031:4]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_ser_in_ready(ram_io_ser_in_ready),
    .io_ser_in_valid(ram_io_ser_in_valid),
    .io_ser_in_bits(ram_io_ser_in_bits),
    .io_ser_out_ready(ram_io_ser_out_ready),
    .io_ser_out_valid(ram_io_ser_out_valid),
    .io_ser_out_bits(ram_io_ser_out_bits),
    .io_tsi_ser_in_ready(ram_io_tsi_ser_in_ready),
    .io_tsi_ser_in_valid(ram_io_tsi_ser_in_valid),
    .io_tsi_ser_in_bits(ram_io_tsi_ser_in_bits),
    .io_tsi_ser_out_ready(ram_io_tsi_ser_out_ready),
    .io_tsi_ser_out_valid(ram_io_tsi_ser_out_valid),
    .io_tsi_ser_out_bits(ram_io_tsi_ser_out_bits)
  );


  SimSerial success_sim ( // @[SerialAdapter.scala 37:23 chipyard.TestHarness.SmallBoomConfig.fir 394041:4]
    .clock(success_sim_clock),
    .reset(success_sim_reset),
    .serial_in_ready(success_sim_serial_in_ready),
    .serial_in_valid(success_sim_serial_in_valid),
    .serial_in_bits(success_sim_serial_in_bits),
    .serial_out_ready(success_sim_serial_out_ready),
    .serial_out_valid(success_sim_serial_out_valid),
    .serial_out_bits(success_sim_serial_out_bits),
    .exit(success_sim_exit)
  );


  SimDRAM #(.LINE_SIZE(64), .ID_BITS(4), .ADDR_BITS(32), .MEM_SIZE(268435456), .DATA_BITS(64)) simdram ( // @[HarnessBinders.scala 146:23 chipyard.TestHarness.SmallBoomConfig.fir 394057:4]
    .clock(simdram_clock),
    .reset(simdram_reset),
    .axi_aw_ready(simdram_axi_aw_ready),
    .axi_aw_valid(simdram_axi_aw_valid),
    .axi_aw_bits_id(simdram_axi_aw_bits_id),
    .axi_aw_bits_addr(simdram_axi_aw_bits_addr),
    .axi_aw_bits_len(simdram_axi_aw_bits_len),
    .axi_aw_bits_size(simdram_axi_aw_bits_size),
    .axi_aw_bits_burst(simdram_axi_aw_bits_burst),
    .axi_aw_bits_lock(simdram_axi_aw_bits_lock),
    .axi_aw_bits_cache(simdram_axi_aw_bits_cache),
    .axi_aw_bits_prot(simdram_axi_aw_bits_prot),
    .axi_aw_bits_qos(simdram_axi_aw_bits_qos),
    .axi_w_ready(simdram_axi_w_ready),
    .axi_w_valid(simdram_axi_w_valid),
    .axi_w_bits_data(simdram_axi_w_bits_data),
    .axi_w_bits_strb(simdram_axi_w_bits_strb),
    .axi_w_bits_last(simdram_axi_w_bits_last),
    .axi_b_ready(simdram_axi_b_ready),
    .axi_b_valid(simdram_axi_b_valid),
    .axi_b_bits_id(simdram_axi_b_bits_id),
    .axi_b_bits_resp(simdram_axi_b_bits_resp),
    .axi_ar_ready(simdram_axi_ar_ready),
    .axi_ar_valid(simdram_axi_ar_valid),
    .axi_ar_bits_id(simdram_axi_ar_bits_id),
    .axi_ar_bits_addr(simdram_axi_ar_bits_addr),
    .axi_ar_bits_len(simdram_axi_ar_bits_len),
    .axi_ar_bits_size(simdram_axi_ar_bits_size),
    .axi_ar_bits_burst(simdram_axi_ar_bits_burst),
    .axi_ar_bits_lock(simdram_axi_ar_bits_lock),
    .axi_ar_bits_cache(simdram_axi_ar_bits_cache),
    .axi_ar_bits_prot(simdram_axi_ar_bits_prot),
    .axi_ar_bits_qos(simdram_axi_ar_bits_qos),
    .axi_r_ready(simdram_axi_r_ready),
    .axi_r_valid(simdram_axi_r_valid),
    .axi_r_bits_id(simdram_axi_r_bits_id),
    .axi_r_bits_data(simdram_axi_r_bits_data),
    .axi_r_bits_resp(simdram_axi_r_bits_resp),
    .axi_r_bits_last(simdram_axi_r_bits_last)
  );


  UARTAdapter_inTestHarness uart_sim_0 ( // @[UARTAdapter.scala 132:28 chipyard.TestHarness.SmallBoomConfig.fir 394064:4]
    .clock(uart_sim_0_clock),
    .reset(uart_sim_0_reset),
    .io_uart_txd(uart_sim_0_io_uart_txd),
    .io_uart_rxd(uart_sim_0_io_uart_rxd)
  );


  assign io_success = success_sim_exit | dtm_success; // @[HarnessBinders.scala 236:22 chipyard.TestHarness.SmallBoomConfig.fir 394054:4 HarnessBinders.scala 236:35 chipyard.TestHarness.SmallBoomConfig.fir 394055:6]
  assign chiptop_jtag_TCK = SimJTAG_jtag_TCK; // @[Periphery.scala 220:15 chipyard.TestHarness.SmallBoomConfig.fir 394004:4]
  assign chiptop_jtag_TMS = SimJTAG_jtag_TMS; // @[Periphery.scala 221:15 chipyard.TestHarness.SmallBoomConfig.fir 394005:4]
  assign chiptop_jtag_TDI = SimJTAG_jtag_TDI; // @[Periphery.scala 222:15 chipyard.TestHarness.SmallBoomConfig.fir 394006:4]
  assign chiptop_serial_tl_bits_in_valid = ram_io_ser_in_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394038:4]
  assign chiptop_serial_tl_bits_in_bits = ram_io_ser_in_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394037:4]
  assign chiptop_serial_tl_bits_out_ready = ram_io_ser_out_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394036:4]
  assign chiptop_axi4_mem_0_bits_aw_ready = simdram_axi_aw_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_w_ready = simdram_axi_w_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_b_valid = simdram_axi_b_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_b_bits_id = simdram_axi_b_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_b_bits_resp = simdram_axi_b_bits_resp; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_ar_ready = simdram_axi_ar_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_r_valid = simdram_axi_r_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_r_bits_id = simdram_axi_r_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_r_bits_data = simdram_axi_r_bits_data; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_r_bits_resp = simdram_axi_r_bits_resp; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_axi4_mem_0_bits_r_bits_last = simdram_axi_r_bits_last; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign chiptop_uart_0_rxd = uart_sim_0_io_uart_rxd; // @[UARTAdapter.scala 135:18 chipyard.TestHarness.SmallBoomConfig.fir 394068:4]
  assign chiptop_reset_wire_reset = reset; // @[TestHarness.scala 41:24 chipyard.TestHarness.SmallBoomConfig.fir 393986:4]
  assign chiptop_clock = clock; // @[Clocks.scala 106:18 chipyard.TestHarness.SmallBoomConfig.fir 393988:4]
  assign SimJTAG_clock = clock; // @[Periphery.scala 225:14 chipyard.TestHarness.SmallBoomConfig.fir 394009:4]
  assign SimJTAG_reset = reset; // @[HarnessBinders.scala 190:97 chipyard.TestHarness.SmallBoomConfig.fir 394001:4]
  assign SimJTAG_jtag_TDO_data = chiptop_jtag_TDO_data; // @[Periphery.scala 223:17 chipyard.TestHarness.SmallBoomConfig.fir 394008:4]
  assign SimJTAG_jtag_TDO_driven = chiptop_jtag_TDO_driven; // @[Periphery.scala 223:17 chipyard.TestHarness.SmallBoomConfig.fir 394007:4]
  assign SimJTAG_enable = plusarg_reader_out[0]; // @[Periphery.scala 228:18 chipyard.TestHarness.SmallBoomConfig.fir 394013:4]
  assign SimJTAG_init_done = ~reset; // @[HarnessBinders.scala 190:105 chipyard.TestHarness.SmallBoomConfig.fir 394003:4]
  assign ram_clock = chiptop_serial_tl_clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 394032:4]
  assign ram_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 393984:4 chipyard.TestHarness.SmallBoomConfig.fir 393985:4]
  assign ram_io_ser_in_ready = chiptop_serial_tl_bits_in_ready; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394039:4]
  assign ram_io_ser_out_valid = chiptop_serial_tl_bits_out_valid; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394035:4]
  assign ram_io_ser_out_bits = chiptop_serial_tl_bits_out_bits; // @[SerialAdapter.scala 28:21 chipyard.TestHarness.SmallBoomConfig.fir 394034:4]
  assign ram_io_tsi_ser_in_valid = success_sim_serial_in_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394052:4]
  assign ram_io_tsi_ser_in_bits = success_sim_serial_in_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394051:4]
  assign ram_io_tsi_ser_out_ready = success_sim_serial_out_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394050:4]
  assign success_sim_clock = chiptop_serial_tl_clock; // @[SerialAdapter.scala 38:20 chipyard.TestHarness.SmallBoomConfig.fir 394046:4]
  assign success_sim_reset = reset; // @[HarnessBinders.scala 235:103 chipyard.TestHarness.SmallBoomConfig.fir 394040:4]
  assign success_sim_serial_in_ready = ram_io_tsi_ser_in_ready; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394053:4]
  assign success_sim_serial_out_valid = ram_io_tsi_ser_out_valid; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394049:4]
  assign success_sim_serial_out_bits = ram_io_tsi_ser_out_bits; // @[SerialAdapter.scala 40:21 chipyard.TestHarness.SmallBoomConfig.fir 394048:4]
  assign simdram_clock = chiptop_axi4_mem_0_clock; // @[HarnessBinders.scala 148:20 chipyard.TestHarness.SmallBoomConfig.fir 394062:4]
  assign simdram_reset = chiptop_axi4_mem_0_reset; // @[HarnessBinders.scala 149:20 chipyard.TestHarness.SmallBoomConfig.fir 394063:4]
  assign simdram_axi_aw_valid = chiptop_axi4_mem_0_bits_aw_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_id = chiptop_axi4_mem_0_bits_aw_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_addr = chiptop_axi4_mem_0_bits_aw_bits_addr; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_len = chiptop_axi4_mem_0_bits_aw_bits_len; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_size = chiptop_axi4_mem_0_bits_aw_bits_size; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_burst = chiptop_axi4_mem_0_bits_aw_bits_burst; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_lock = chiptop_axi4_mem_0_bits_aw_bits_lock; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_cache = chiptop_axi4_mem_0_bits_aw_bits_cache; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_prot = chiptop_axi4_mem_0_bits_aw_bits_prot; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_aw_bits_qos = chiptop_axi4_mem_0_bits_aw_bits_qos; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_w_valid = chiptop_axi4_mem_0_bits_w_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_w_bits_data = chiptop_axi4_mem_0_bits_w_bits_data; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_w_bits_strb = chiptop_axi4_mem_0_bits_w_bits_strb; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_w_bits_last = chiptop_axi4_mem_0_bits_w_bits_last; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_b_ready = chiptop_axi4_mem_0_bits_b_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_valid = chiptop_axi4_mem_0_bits_ar_valid; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_id = chiptop_axi4_mem_0_bits_ar_bits_id; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_addr = chiptop_axi4_mem_0_bits_ar_bits_addr; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_len = chiptop_axi4_mem_0_bits_ar_bits_len; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_size = chiptop_axi4_mem_0_bits_ar_bits_size; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_burst = chiptop_axi4_mem_0_bits_ar_bits_burst; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_lock = chiptop_axi4_mem_0_bits_ar_bits_lock; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_cache = chiptop_axi4_mem_0_bits_ar_bits_cache; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_prot = chiptop_axi4_mem_0_bits_ar_bits_prot; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_ar_bits_qos = chiptop_axi4_mem_0_bits_ar_bits_qos; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign simdram_axi_r_ready = chiptop_axi4_mem_0_bits_r_ready; // @[HarnessBinders.scala 147:18 chipyard.TestHarness.SmallBoomConfig.fir 394061:4]
  assign uart_sim_0_clock = clock; // @[chipyard.TestHarness.SmallBoomConfig.fir 394065:4]
  assign uart_sim_0_reset = reset; // @[chipyard.TestHarness.SmallBoomConfig.fir 394066:4]
  assign uart_sim_0_io_uart_txd = chiptop_uart_0_txd; // @[UARTAdapter.scala 134:28 chipyard.TestHarness.SmallBoomConfig.fir 394067:4]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fwrite(32'h80000002,"*** FAILED *** (exit code = %d)\n",_T_4); // @[Periphery.scala 235:13 chipyard.TestHarness.SmallBoomConfig.fir 394023:8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3 & _T_2) begin
          $fatal; // @[Periphery.scala 236:11 chipyard.TestHarness.SmallBoomConfig.fir 394028:8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule



module mem_inTestHarness(
  input  [8:0] RW0_addr,
  input        RW0_en,
  input        RW0_clk,
  input        RW0_wmode,
  input  [7:0] RW0_wdata_0,
  input  [7:0] RW0_wdata_1,
  input  [7:0] RW0_wdata_2,
  input  [7:0] RW0_wdata_3,
  input  [7:0] RW0_wdata_4,
  input  [7:0] RW0_wdata_5,
  input  [7:0] RW0_wdata_6,
  input  [7:0] RW0_wdata_7,
  output [7:0] RW0_rdata_0,
  output [7:0] RW0_rdata_1,
  output [7:0] RW0_rdata_2,
  output [7:0] RW0_rdata_3,
  output [7:0] RW0_rdata_4,
  output [7:0] RW0_rdata_5,
  output [7:0] RW0_rdata_6,
  output [7:0] RW0_rdata_7,
  input        RW0_wmask_0,
  input        RW0_wmask_1,
  input        RW0_wmask_2,
  input        RW0_wmask_3,
  input        RW0_wmask_4,
  input        RW0_wmask_5,
  input        RW0_wmask_6,
  input        RW0_wmask_7
);
  wire [8:0] mem_ext_RW0_addr;
  wire  mem_ext_RW0_en;
  wire  mem_ext_RW0_clk;
  wire  mem_ext_RW0_wmode;
  wire [63:0] mem_ext_RW0_wdata;
  wire [63:0] mem_ext_RW0_rdata;
  wire [7:0] mem_ext_RW0_wmask;
  wire [31:0] _GEN_4 = {RW0_wdata_7,RW0_wdata_6,RW0_wdata_5,RW0_wdata_4};
  wire [31:0] _GEN_5 = {RW0_wdata_3,RW0_wdata_2,RW0_wdata_1,RW0_wdata_0};
  wire [3:0] _GEN_10 = {RW0_wmask_7,RW0_wmask_6,RW0_wmask_5,RW0_wmask_4};
  wire [3:0] _GEN_11 = {RW0_wmask_3,RW0_wmask_2,RW0_wmask_1,RW0_wmask_0};
  mem_ext mem_ext (
    .RW0_addr(mem_ext_RW0_addr),
    .RW0_en(mem_ext_RW0_en),
    .RW0_clk(mem_ext_RW0_clk),
    .RW0_wmode(mem_ext_RW0_wmode),
    .RW0_wdata(mem_ext_RW0_wdata),
    .RW0_rdata(mem_ext_RW0_rdata),
    .RW0_wmask(mem_ext_RW0_wmask)
  );
  assign mem_ext_RW0_clk = RW0_clk;
  assign mem_ext_RW0_en = RW0_en;
  assign mem_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = mem_ext_RW0_rdata[7:0];
  assign RW0_rdata_1 = mem_ext_RW0_rdata[15:8];
  assign RW0_rdata_2 = mem_ext_RW0_rdata[23:16];
  assign RW0_rdata_3 = mem_ext_RW0_rdata[31:24];
  assign RW0_rdata_4 = mem_ext_RW0_rdata[39:32];
  assign RW0_rdata_5 = mem_ext_RW0_rdata[47:40];
  assign RW0_rdata_6 = mem_ext_RW0_rdata[55:48];
  assign RW0_rdata_7 = mem_ext_RW0_rdata[63:56];
  assign mem_ext_RW0_wmode = RW0_wmode;
  assign mem_ext_RW0_wdata = {_GEN_4,_GEN_5};
  assign mem_ext_RW0_wmask = {_GEN_10,_GEN_11};
endmodule
